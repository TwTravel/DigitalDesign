// Implements a simple Nios II system for the DE2 board.
// Inputs: SW7-0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7-0 are parallel port outputs from the Nios II system
module TimerTest(SW, KEY, CLOCK_50, LEDG, HEX7, HEX6, HEX5, HEX4);
input [7:0] SW;
input [0:0] KEY;
input CLOCK_50;
output [7:0] LEDG;
output [6:0] HEX6, HEX7, HEX5, HEX4;
// Instantiate the Nios II system module generated by the SOPC Builder:
// nios_system (clk, reset_n, out_port_from_the_LEDs, in_port_to_the_Switches)
NiosII niosIItimer(CLOCK_50, KEY[0], LEDG, SW);

//output switch settings
HexDigit Digit7(HEX7, SW[7:4]);
HexDigit Digit6(HEX6, SW[3:0]);
//output LEDs
HexDigit Digit5(HEX5, LEDG[7:4]);
HexDigit Digit4(HEX4, LEDG[3:0]);


endmodule

//////////////////////////////////////////////
// Decode one hex digit for LED 7-seg display
module HexDigit(segs, num);
	input [3:0] num	;		//the hex digit to be displayed
	output [6:0] segs ;		//actual LED segments
	reg [6:0] segs ;
	always @ (num)
	begin
		case (num)
				4'h0: segs = 7'b1000000;
				4'h1: segs = 7'b1111001;
				4'h2: segs = 7'b0100100;
				4'h3: segs = 7'b0110000;
				4'h4: segs = 7'b0011001;
				4'h5: segs = 7'b0010010;
				4'h6: segs = 7'b0000010;
				4'h7: segs = 7'b1111000;
				4'h8: segs = 7'b0000000;
				4'h9: segs = 7'b0010000;
				4'ha: segs = 7'b0001000;
				4'hb: segs = 7'b0000011;
				4'hc: segs = 7'b1000110;
				4'hd: segs = 7'b0100001;
				4'he: segs = 7'b0000110;
				4'hf: segs = 7'b0001110;
				default segs = 7'b1111111;
		endcase
	end
endmodule
///////////////////////////////////////////////