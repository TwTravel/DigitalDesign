// Implements a  Nios II system with SDRAM and DDS control for the DE2 board.
// Inputs: SW7-0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7-0 are parallel port outputs from the Nios II system
module TimerSDRAM(SW, KEY, CLOCK_50, LEDG, 
	HEX3, HEX2, HEX1, HEX0, HEX5, HEX4, 
	GPIO_0,
	DRAM_CLK, DRAM_CKE,
	DRAM_ADDR, DRAM_BA_1, DRAM_BA_0, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,
	DRAM_WE_N, DRAM_DQ, DRAM_UDQM, DRAM_LDQM,
	VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_R, VGA_G, VGA_B  
	);
	
	input [15:0] SW;
	input [0:0] KEY;
	input CLOCK_50;
	output [7:0] LEDG;
	output [6:0] HEX3, HEX2, HEX1, HEX0, HEX5, HEX4;
	output [35:0] GPIO_0;
	//SDRAM
	output [11:0] DRAM_ADDR;
	output DRAM_BA_1, DRAM_BA_0, DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK;
	output DRAM_CKE, DRAM_CS_N, DRAM_WE_N, DRAM_UDQM, DRAM_LDQM;
	inout [15:0] DRAM_DQ;
	//VGA
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK;				//	VGA BLANK
	output			VGA_SYNC;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	
	reg [31:0] DDS_accum;
	wire [31:0] DDS_incr;
	
	// Instantiate the Nios II system module generated by the SOPC Builder:
	//module NiosSDRAM (clk, reset_n, out_port_from_the_LED,
	//
    //                zs_addr_from_the_sdram_0,
    //                zs_ba_from_the_sdram_0,
    //                zs_cas_n_from_the_sdram_0,
    //                zs_cke_from_the_sdram_0,
    //                zs_cs_n_from_the_sdram_0,
    //                zs_dq_to_and_from_the_sdram_0,
    //                zs_dqm_from_the_sdram_0,
    //                zs_ras_n_from_the_sdram_0,
    //                zs_we_n_from_the_sdram_0,
    //
    //				  in_port_to_the_switch, out_port_from_the_wideOut )
	NiosSDRAM nios2(CLOCK_50, KEY[0], LEDG, 
				DRAM_ADDR,
				{DRAM_BA_1, DRAM_BA_0},
				DRAM_CAS_N,
				DRAM_CKE,
				DRAM_CS_N,
				DRAM_DQ,
				{DRAM_UDQM, DRAM_LDQM},
				DRAM_RAS_N,
				DRAM_WE_N,
				SW[7:0], DDS_incr);
				
	// Instantiate the module sdram_pll (inclk0, c0)
	// to shift sdram clock -3 ns as suggested in
	// tut_DE2_sdram_verilog.pdf
	sdram_pll neg_3ns (CLOCK_50, DRAM_CLK);

	//show switch settings
	HexDigit Digit3(HEX3, SW[15:12]);
	HexDigit Digit2(HEX2, SW[11:8]);
	HexDigit Digit1(HEX1, SW[7:4]);
	HexDigit Digit0(HEX0, SW[3:0]);
	//show LEDs as hex
	HexDigit Digit5(HEX5, LEDG[7:4]);
	HexDigit Digit4(HEX4, LEDG[3:0]);
	
	//make a direct digital systnesis accumulator 
	// and output the top 8 bits
	always @ (posedge CLOCK_50) begin
		DDS_accum <= DDS_accum + DDS_incr ;
	end
	assign GPIO_0[7:0] = DDS_accum[31:24];
	//use the VGA DAC for an audio signal 
	assign VGA_R =  DDS_accum[31:22]; //10-bits
	assign VGA_SYNC = 1;
	assign VGA_BLANK = 1;
	assign VGA_CLK = CLOCK_50;
	
endmodule

//////////////////////////////////////////////
// Decode one hex digit for LED 7-seg display
module HexDigit(segs, num);
	input [3:0] num	;		//the hex digit to be displayed
	output [6:0] segs ;		//actual LED segments
	reg [6:0] segs ;
	always @ (num)
	begin
		case (num)
				4'h0: segs = 7'b1000000;
				4'h1: segs = 7'b1111001;
				4'h2: segs = 7'b0100100;
				4'h3: segs = 7'b0110000;
				4'h4: segs = 7'b0011001;
				4'h5: segs = 7'b0010010;
				4'h6: segs = 7'b0000010;
				4'h7: segs = 7'b1111000;
				4'h8: segs = 7'b0000000;
				4'h9: segs = 7'b0010000;
				4'ha: segs = 7'b0001000;
				4'hb: segs = 7'b0000011;
				4'hc: segs = 7'b1000110;
				4'hd: segs = 7'b0100001;
				4'he: segs = 7'b0000110;
				4'hf: segs = 7'b0001110;
				default segs = 7'b1111111;
		endcase
	end
endmodule
///////////////////////////////////////////////