// Implements a  Nios II system with SDRAM and DDS control for the DE2 board.
// Inputs: SW7-0 are parallel port inputs to the Nios II system
// CLOCK_50 is the system clock
// KEY0 is the active-low system reset
// Outputs: LEDG7-0 are parallel port outputs from the Nios II system
module TestBigNios(SW, KEY, CLOCK_50, LEDG, 
	HEX3, HEX2, HEX1, HEX0, HEX5, HEX4, 
	GPIO_0,
	DRAM_CLK, DRAM_CKE,
	DRAM_ADDR, DRAM_BA_1, DRAM_BA_0, DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N,
	DRAM_WE_N, DRAM_DQ, DRAM_UDQM, DRAM_LDQM,
	VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_R, VGA_G, VGA_B,
	LCD_ON, LCD_BLON, LCD_RW, LCD_EN, LCD_RS, LCD_DATA				  
	);
	
	input [17:0] SW;
	input [3:0] KEY;
	input CLOCK_50;
	output [7:0] LEDG;
	output [6:0] HEX3, HEX2, HEX1, HEX0, HEX5, HEX4;
	output [35:0] GPIO_0;
	//SDRAM
	output [11:0] DRAM_ADDR;
	output DRAM_BA_1, DRAM_BA_0, DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK;
	output DRAM_CKE, DRAM_CS_N, DRAM_WE_N, DRAM_UDQM, DRAM_LDQM;
	inout [15:0] DRAM_DQ;
	//VGA
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK;				//	VGA BLANK
	output			VGA_SYNC;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	//LCD
	inout	[7:0]	LCD_DATA;				//	LCD Data bus 8 bits
	output			LCD_ON;					//	LCD Power ON/OFF
	output			LCD_BLON;				//	LCD Back Light ON/OFF
	output			LCD_RW;					//	LCD Read/Write Select, 0 = Write, 1 = Read
	output			LCD_EN;					//	LCD Enable
	output			LCD_RS;					//	LCD Command/Data Select, 0 = Command, 1 = Data  
	
	//DDS hardware
	reg [31:0] DDS_accum;
	wire [31:0] DDS_incr, Out1;
	wire [9:0] sine_out, cos_out;
	
	// Instantiate the Nios II system module generated by the SOPC Builder:
	//from the file bigNios.v
	//module bigNios (clk, reset_n,
	//				in_port_to_the_In0, 
	//				in_port_to_the_In1_8bit,
	//				out_port_from_the_Out0, 
	//				out_port_from_the_Out1,
    //           // the_lcd
    //             LCD_E_from_the_lcd,
    //              LCD_RS_from_the_lcd,
    //              LCD_RW_from_the_lcd,
    //              LCD_data_to_and_from_the_lcd,
    //           // the_sdram_0
    //              zs_addr_from_the_sdram_0,
    //              zs_ba_from_the_sdram_0,
    //              zs_cas_n_from_the_sdram_0,
    //              zs_cke_from_the_sdram_0,
    //              zs_cs_n_from_the_sdram_0,
    //              zs_dq_to_and_from_the_sdram_0,
    //              zs_dqm_from_the_sdram_0,
    //              zs_ras_n_from_the_sdram_0,
    //              zs_we_n_from_the_sdram_0  )

	bigNios nios2(CLOCK_50, KEY[0],
				// parallel i/o
				SW,			//In0 32 bits
				KEY,		//In1 8 bits
				DDS_incr,	//Out0
				Out1,		//Out1
				// lcd
				LCD_EN, LCD_RS, LCD_RW, LCD_DATA,
        		// sdram 
				DRAM_ADDR,
				{DRAM_BA_1, DRAM_BA_0},
				DRAM_CAS_N,
				DRAM_CKE,
				DRAM_CS_N,
				DRAM_DQ,
				{DRAM_UDQM, DRAM_LDQM},
				DRAM_RAS_N,
				DRAM_WE_N);
				
	// Instantiate the module sdram_pll (inclk0, c0)
	// to shift sdram clock -3 ns as suggested in
	// tut_DE2_sdram_verilog.pdf
	sdram_pll neg_3ns (CLOCK_50, DRAM_CLK);

	//show switch settings
	HexDigit Digit3(HEX3, SW[15:12]);
	HexDigit Digit2(HEX2, SW[11:8]);
	HexDigit Digit1(HEX1, SW[7:4]);
	HexDigit Digit0(HEX0, SW[3:0]);
	//show LEDs as hex
	HexDigit Digit5(HEX5, LEDG[7:4]);
	HexDigit Digit4(HEX4, LEDG[3:0]);
	
	//make a direct digital systnesis accumulator 
	// and output the top 8 bits to connector JP1
	// and output a 10-bit sine wave to the VGA plug
	always @ (posedge CLOCK_50) begin
		DDS_accum <= DDS_accum + DDS_incr ;
	end
	assign GPIO_0[7:0] = DDS_accum[31:24];
	
	//hook up the ROM table
	sync_rom sineTable(CLOCK_50, DDS_accum[31:24], sine_out);
	sync_rom cosTable(CLOCK_50, DDS_accum[31:24]+8'h40, cos_out);
	
	//use the VGA DAC for an audio signal 
	assign VGA_R = sine_out ; //10-bits
	assign VGA_B = cos_out ; //10-bits
	assign VGA_SYNC = 1 ;
	assign VGA_BLANK = 1 ;
	assign VGA_CLK = CLOCK_50 ;
	
	//disable the LCD for now
	assign LCD_ON = 0;
	assign LCD_BLON = 0;
	
endmodule

//////////////////////////////////////////////
// Decode one hex digit for LED 7-seg display
module HexDigit(segs, num);
	input [3:0] num	;		//the hex digit to be displayed
	output [6:0] segs ;		//actual LED segments
	reg [6:0] segs ;
	always @ (num)
	begin
		case (num)
				4'h0: segs = 7'b1000000;
				4'h1: segs = 7'b1111001;
				4'h2: segs = 7'b0100100;
				4'h3: segs = 7'b0110000;
				4'h4: segs = 7'b0011001;
				4'h5: segs = 7'b0010010;
				4'h6: segs = 7'b0000010;
				4'h7: segs = 7'b1111000;
				4'h8: segs = 7'b0000000;
				4'h9: segs = 7'b0010000;
				4'ha: segs = 7'b0001000;
				4'hb: segs = 7'b0000011;
				4'hc: segs = 7'b1000110;
				4'hd: segs = 7'b0100001;
				4'he: segs = 7'b0000110;
				4'hf: segs = 7'b0001110;
				default segs = 7'b1111111;
		endcase
	end
endmodule
///////////////////////////////////////////////
// Infer ROM storage
// for a sin table for the DDS

module sync_rom (clock, address, sine);
	input clock;
	input [7:0] address;
	output [9:0] sine;
	reg [9:0] sine;
	always @ (posedge clock)
	begin
		case (address)
			8'h00: sine = 10'h200 ;
			8'h01: sine = 10'h20c ;
			8'h02: sine = 10'h219 ;
			8'h03: sine = 10'h225 ;
			8'h04: sine = 10'h232 ;
			8'h05: sine = 10'h23e ;
			8'h06: sine = 10'h24a ;
			8'h07: sine = 10'h257 ;
			8'h08: sine = 10'h263 ;
			8'h09: sine = 10'h26f ;
			8'h0a: sine = 10'h27c ;
			8'h0b: sine = 10'h288 ;
			8'h0c: sine = 10'h294 ;
			8'h0d: sine = 10'h2a0 ;
			8'h0e: sine = 10'h2ac ;
			8'h0f: sine = 10'h2b7 ;
			8'h10: sine = 10'h2c3 ;
			8'h11: sine = 10'h2cf ;
			8'h12: sine = 10'h2da ;
			8'h13: sine = 10'h2e5 ;
			8'h14: sine = 10'h2f0 ;
			8'h15: sine = 10'h2fb ;
			8'h16: sine = 10'h306 ;
			8'h17: sine = 10'h311 ;
			8'h18: sine = 10'h31b ;
			8'h19: sine = 10'h326 ;
			8'h1a: sine = 10'h330 ;
			8'h1b: sine = 10'h33a ;
			8'h1c: sine = 10'h344 ;
			8'h1d: sine = 10'h34d ;
			8'h1e: sine = 10'h357 ;
			8'h1f: sine = 10'h360 ;
			8'h20: sine = 10'h369 ;
			8'h21: sine = 10'h372 ;
			8'h22: sine = 10'h37a ;
			8'h23: sine = 10'h382 ;
			8'h24: sine = 10'h38b ;
			8'h25: sine = 10'h392 ;
			8'h26: sine = 10'h39a ;
			8'h27: sine = 10'h3a1 ;
			8'h28: sine = 10'h3a8 ;
			8'h29: sine = 10'h3af ;
			8'h2a: sine = 10'h3b6 ;
			8'h2b: sine = 10'h3bc ;
			8'h2c: sine = 10'h3c2 ;
			8'h2d: sine = 10'h3c8 ;
			8'h2e: sine = 10'h3cd ;
			8'h2f: sine = 10'h3d3 ;
			8'h30: sine = 10'h3d8 ;
			8'h31: sine = 10'h3dc ;
			8'h32: sine = 10'h3e1 ;
			8'h33: sine = 10'h3e5 ;
			8'h34: sine = 10'h3e8 ;
			8'h35: sine = 10'h3ec ;
			8'h36: sine = 10'h3ef ;
			8'h37: sine = 10'h3f2 ;
			8'h38: sine = 10'h3f5 ;
			8'h39: sine = 10'h3f7 ;
			8'h3a: sine = 10'h3f9 ;
			8'h3b: sine = 10'h3fb ;
			8'h3c: sine = 10'h3fc ;
			8'h3d: sine = 10'h3fd ;
			8'h3e: sine = 10'h3fe ;
			8'h3f: sine = 10'h3fe ;
			8'h40: sine = 10'h3ff ;
			8'h41: sine = 10'h3fe ;
			8'h42: sine = 10'h3fe ;
			8'h43: sine = 10'h3fd ;
			8'h44: sine = 10'h3fc ;
			8'h45: sine = 10'h3fb ;
			8'h46: sine = 10'h3f9 ;
			8'h47: sine = 10'h3f7 ;
			8'h48: sine = 10'h3f5 ;
			8'h49: sine = 10'h3f2 ;
			8'h4a: sine = 10'h3ef ;
			8'h4b: sine = 10'h3ec ;
			8'h4c: sine = 10'h3e8 ;
			8'h4d: sine = 10'h3e5 ;
			8'h4e: sine = 10'h3e1 ;
			8'h4f: sine = 10'h3dc ;
			8'h50: sine = 10'h3d8 ;
			8'h51: sine = 10'h3d3 ;
			8'h52: sine = 10'h3cd ;
			8'h53: sine = 10'h3c8 ;
			8'h54: sine = 10'h3c2 ;
			8'h55: sine = 10'h3bc ;
			8'h56: sine = 10'h3b6 ;
			8'h57: sine = 10'h3af ;
			8'h58: sine = 10'h3a8 ;
			8'h59: sine = 10'h3a1 ;
			8'h5a: sine = 10'h39a ;
			8'h5b: sine = 10'h392 ;
			8'h5c: sine = 10'h38b ;
			8'h5d: sine = 10'h382 ;
			8'h5e: sine = 10'h37a ;
			8'h5f: sine = 10'h372 ;
			8'h60: sine = 10'h369 ;
			8'h61: sine = 10'h360 ;
			8'h62: sine = 10'h357 ;
			8'h63: sine = 10'h34d ;
			8'h64: sine = 10'h344 ;
			8'h65: sine = 10'h33a ;
			8'h66: sine = 10'h330 ;
			8'h67: sine = 10'h326 ;
			8'h68: sine = 10'h31b ;
			8'h69: sine = 10'h311 ;
			8'h6a: sine = 10'h306 ;
			8'h6b: sine = 10'h2fb ;
			8'h6c: sine = 10'h2f0 ;
			8'h6d: sine = 10'h2e5 ;
			8'h6e: sine = 10'h2da ;
			8'h6f: sine = 10'h2cf ;
			8'h70: sine = 10'h2c3 ;
			8'h71: sine = 10'h2b7 ;
			8'h72: sine = 10'h2ac ;
			8'h73: sine = 10'h2a0 ;
			8'h74: sine = 10'h294 ;
			8'h75: sine = 10'h288 ;
			8'h76: sine = 10'h27c ;
			8'h77: sine = 10'h26f ;
			8'h78: sine = 10'h263 ;
			8'h79: sine = 10'h257 ;
			8'h7a: sine = 10'h24a ;
			8'h7b: sine = 10'h23e ;
			8'h7c: sine = 10'h232 ;
			8'h7d: sine = 10'h225 ;
			8'h7e: sine = 10'h219 ;
			8'h7f: sine = 10'h20c ;
			8'h80: sine = 10'h200 ;
			8'h81: sine = 10'h1f3 ;
			8'h82: sine = 10'h1e6 ;
			8'h83: sine = 10'h1da ;
			8'h84: sine = 10'h1cd ;
			8'h85: sine = 10'h1c1 ;
			8'h86: sine = 10'h1b5 ;
			8'h87: sine = 10'h1a8 ;
			8'h88: sine = 10'h19c ;
			8'h89: sine = 10'h190 ;
			8'h8a: sine = 10'h183 ;
			8'h8b: sine = 10'h177 ;
			8'h8c: sine = 10'h16b ;
			8'h8d: sine = 10'h15f ;
			8'h8e: sine = 10'h153 ;
			8'h8f: sine = 10'h148 ;
			8'h90: sine = 10'h13c ;
			8'h91: sine = 10'h130 ;
			8'h92: sine = 10'h125 ;
			8'h93: sine = 10'h11a ;
			8'h94: sine = 10'h10f ;
			8'h95: sine = 10'h104 ;
			8'h96: sine = 10'h0f9 ;
			8'h97: sine = 10'h0ee ;
			8'h98: sine = 10'h0e4 ;
			8'h99: sine = 10'h0d9 ;
			8'h9a: sine = 10'h0cf ;
			8'h9b: sine = 10'h0c5 ;
			8'h9c: sine = 10'h0bb ;
			8'h9d: sine = 10'h0b2 ;
			8'h9e: sine = 10'h0a8 ;
			8'h9f: sine = 10'h09f ;
			8'ha0: sine = 10'h096 ;
			8'ha1: sine = 10'h08d ;
			8'ha2: sine = 10'h085 ;
			8'ha3: sine = 10'h07d ;
			8'ha4: sine = 10'h074 ;
			8'ha5: sine = 10'h06d ;
			8'ha6: sine = 10'h065 ;
			8'ha7: sine = 10'h05e ;
			8'ha8: sine = 10'h057 ;
			8'ha9: sine = 10'h050 ;
			8'haa: sine = 10'h049 ;
			8'hab: sine = 10'h043 ;
			8'hac: sine = 10'h03d ;
			8'had: sine = 10'h037 ;
			8'hae: sine = 10'h032 ;
			8'haf: sine = 10'h02c ;
			8'hb0: sine = 10'h027 ;
			8'hb1: sine = 10'h023 ;
			8'hb2: sine = 10'h01e ;
			8'hb3: sine = 10'h01a ;
			8'hb4: sine = 10'h017 ;
			8'hb5: sine = 10'h013 ;
			8'hb6: sine = 10'h010 ;
			8'hb7: sine = 10'h00d ;
			8'hb8: sine = 10'h00a ;
			8'hb9: sine = 10'h008 ;
			8'hba: sine = 10'h006 ;
			8'hbb: sine = 10'h004 ;
			8'hbc: sine = 10'h003 ;
			8'hbd: sine = 10'h002 ;
			8'hbe: sine = 10'h001 ;
			8'hbf: sine = 10'h001 ;
			8'hc0: sine = 10'h001 ;
			8'hc1: sine = 10'h001 ;
			8'hc2: sine = 10'h001 ;
			8'hc3: sine = 10'h002 ;
			8'hc4: sine = 10'h003 ;
			8'hc5: sine = 10'h004 ;
			8'hc6: sine = 10'h006 ;
			8'hc7: sine = 10'h008 ;
			8'hc8: sine = 10'h00a ;
			8'hc9: sine = 10'h00d ;
			8'hca: sine = 10'h010 ;
			8'hcb: sine = 10'h013 ;
			8'hcc: sine = 10'h017 ;
			8'hcd: sine = 10'h01a ;
			8'hce: sine = 10'h01e ;
			8'hcf: sine = 10'h023 ;
			8'hd0: sine = 10'h027 ;
			8'hd1: sine = 10'h02c ;
			8'hd2: sine = 10'h032 ;
			8'hd3: sine = 10'h037 ;
			8'hd4: sine = 10'h03d ;
			8'hd5: sine = 10'h043 ;
			8'hd6: sine = 10'h049 ;
			8'hd7: sine = 10'h050 ;
			8'hd8: sine = 10'h057 ;
			8'hd9: sine = 10'h05e ;
			8'hda: sine = 10'h065 ;
			8'hdb: sine = 10'h06d ;
			8'hdc: sine = 10'h074 ;
			8'hdd: sine = 10'h07d ;
			8'hde: sine = 10'h085 ;
			8'hdf: sine = 10'h08d ;
			8'he0: sine = 10'h096 ;
			8'he1: sine = 10'h09f ;
			8'he2: sine = 10'h0a8 ;
			8'he3: sine = 10'h0b2 ;
			8'he4: sine = 10'h0bb ;
			8'he5: sine = 10'h0c5 ;
			8'he6: sine = 10'h0cf ;
			8'he7: sine = 10'h0d9 ;
			8'he8: sine = 10'h0e4 ;
			8'he9: sine = 10'h0ee ;
			8'hea: sine = 10'h0f9 ;
			8'heb: sine = 10'h104 ;
			8'hec: sine = 10'h10f ;
			8'hed: sine = 10'h11a ;
			8'hee: sine = 10'h125 ;
			8'hef: sine = 10'h130 ;
			8'hf0: sine = 10'h13c ;
			8'hf1: sine = 10'h148 ;
			8'hf2: sine = 10'h153 ;
			8'hf3: sine = 10'h15f ;
			8'hf4: sine = 10'h16b ;
			8'hf5: sine = 10'h177 ;
			8'hf6: sine = 10'h183 ;
			8'hf7: sine = 10'h190 ;
			8'hf8: sine = 10'h19c ;
			8'hf9: sine = 10'h1a8 ;
			8'hfa: sine = 10'h1b5 ;
			8'hfb: sine = 10'h1c1 ;
			8'hfc: sine = 10'h1cd ;
			8'hfd: sine = 10'h1da ;
			8'hfe: sine = 10'h1e6 ;
			8'hff: sine = 10'h1f3 ;
		endcase
	end
endmodule
///////////////////////////////////////////////