// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsqrt 

// ============================================================
// File Name: stage4sqrt.v
// Megafunction Name(s):
// 			altsqrt
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.0 Build 178 04/27/2006 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt2stage (
	clk,
	radical,
	q,
	remainder);
	
parameter BusWidth = 0;
parameter DecimalWidth = 0;

	input	  clk;
	input	[BusWidth*2-1:0]  radical;
	output	[BusWidth-1:0]  q;
	output	[BusWidth:0]  remainder;

	wire [BusWidth:0] sub_wire0;
	wire [BusWidth-1:0] sub_wire1;
	wire [BusWidth:0] remainder = sub_wire0[BusWidth:0];
	wire [BusWidth-1:0] q = sub_wire1[BusWidth-1:0];

	altsqrt	altsqrt_component (
				.radical (radical),
				.clk (clk),
				.remainder (sub_wire0),
				.q (sub_wire1)
				// synopsys translate_off
				,
				.aclr (),
				.ena ()
				// synopsys translate_on
				);
	defparam
		altsqrt_component.pipeline = 2,
		altsqrt_component.q_port_width = BusWidth,
		altsqrt_component.r_port_width = BusWidth+1,
		altsqrt_component.width = BusWidth*2;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "12"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "13"
// Retrieval info: CONSTANT: WIDTH NUMERIC "24"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL clk
// Retrieval info: USED_PORT: q 0 0 12 0 OUTPUT NODEFVAL q[11..0]
// Retrieval info: USED_PORT: radical 0 0 24 0 INPUT NODEFVAL radical[23..0]
// Retrieval info: USED_PORT: remainder 0 0 13 0 OUTPUT NODEFVAL remainder[12..0]
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 24 0 radical 0 0 24 0
// Retrieval info: CONNECT: q 0 0 12 0 @q 0 0 12 0
// Retrieval info: CONNECT: remainder 0 0 13 0 @remainder 0 0 13 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL stage4sqrt_bb.v FALSE
