////////////////////////////////
// Conversion from RGB[10,10,10] to RGB[10,10,10]
// Simplifies Hues, as well as Saturation and Lightness via a look up table
// ECE 5760 - Cornell University - Fall 2010
// Kerran Flanagan, Tom Gowing, Jeff Yates
////////////////////////////////

module RGB_HueSimplifier (
	clock,
	iRed,
	iGreen,
	iBlue,
	oRed,
	oGreen,
	oBlue
	);
	
	input	wire	clock;
	input	wire	unsigned [9:0]	iRed, iGreen, iBlue;
	output 	wire 	unsigned [9:0] 	oRed, oGreen, oBlue;
	
	//use a 3 bit per color lookup table
	
	wire unsigned [2:0] iR, iG, iB;
	
	assign iR = iRed[9:7];
	assign iG = iGreen[9:7];
	assign iB = iBlue[9:7];
	

	wire unsigned [8:0] tableInput;
	
	assign tableInput = {iR, iG, iB};
	
	reg unsigned [8:0] tableResult;
	
	wire unsigned [2:0] oR, oG, oB;
	
	assign oR = tableResult[8:6];
	assign oG = tableResult[5:3];
	assign oB = tableResult[2:0];
	
	assign oRed = {oR,7'd0};
	assign oGreen = {oG,7'd0};
	assign oBlue = {oB,7'd0};
	
	always @(posedge clock) begin
		case (tableInput)
			//begin code from matlab
9'b000000000: tableResult <= {9'b010010010};
9'b000000001: tableResult <= {9'b000000100};
9'b000000010: tableResult <= {9'b000000100};
9'b000000011: tableResult <= {9'b000000100};
9'b000000100: tableResult <= {9'b000000100};
9'b000000101: tableResult <= {9'b000000100};
9'b000000110: tableResult <= {9'b010010111};
9'b000000111: tableResult <= {9'b010010111};
9'b000001000: tableResult <= {9'b000100000};
9'b000001001: tableResult <= {9'b000100100};
9'b000001010: tableResult <= {9'b000010100};
9'b000001011: tableResult <= {9'b000001100};
9'b000001100: tableResult <= {9'b000001100};
9'b000001101: tableResult <= {9'b000001100};
9'b000001110: tableResult <= {9'b010011111};
9'b000001111: tableResult <= {9'b010010111};
9'b000010000: tableResult <= {9'b000100000};
9'b000010001: tableResult <= {9'b000100010};
9'b000010010: tableResult <= {9'b000100100};
9'b000010011: tableResult <= {9'b000010100};
9'b000010100: tableResult <= {9'b000010100};
9'b000010101: tableResult <= {9'b000010100};
9'b000010110: tableResult <= {9'b010011111};
9'b000010111: tableResult <= {9'b010011111};
9'b000011000: tableResult <= {9'b000100000};
9'b000011001: tableResult <= {9'b000100001};
9'b000011010: tableResult <= {9'b000100010};
9'b000011011: tableResult <= {9'b000100100};
9'b000011100: tableResult <= {9'b000011100};
9'b000011101: tableResult <= {9'b000010100};
9'b000011110: tableResult <= {9'b010100111};
9'b000011111: tableResult <= {9'b010100111};
9'b000100000: tableResult <= {9'b000100000};
9'b000100001: tableResult <= {9'b000100001};
9'b000100010: tableResult <= {9'b000100010};
9'b000100011: tableResult <= {9'b000100011};
9'b000100100: tableResult <= {9'b000100100};
9'b000100101: tableResult <= {9'b000011100};
9'b000100110: tableResult <= {9'b010101111};
9'b000100111: tableResult <= {9'b010101111};
9'b000101000: tableResult <= {9'b000100000};
9'b000101001: tableResult <= {9'b000100001};
9'b000101010: tableResult <= {9'b000100010};
9'b000101011: tableResult <= {9'b000100010};
9'b000101100: tableResult <= {9'b000100011};
9'b000101101: tableResult <= {9'b000100100};
9'b000101110: tableResult <= {9'b010110111};
9'b000101111: tableResult <= {9'b010101111};
9'b000110000: tableResult <= {9'b010111010};
9'b000110001: tableResult <= {9'b010111011};
9'b000110010: tableResult <= {9'b010111011};
9'b000110011: tableResult <= {9'b010111100};
9'b000110100: tableResult <= {9'b010111101};
9'b000110101: tableResult <= {9'b010111110};
9'b000110110: tableResult <= {9'b010111111};
9'b000110111: tableResult <= {9'b010110111};
9'b000111000: tableResult <= {9'b010111010};
9'b000111001: tableResult <= {9'b010111010};
9'b000111010: tableResult <= {9'b010111011};
9'b000111011: tableResult <= {9'b010111100};
9'b000111100: tableResult <= {9'b010111101};
9'b000111101: tableResult <= {9'b010111101};
9'b000111110: tableResult <= {9'b010111110};
9'b000111111: tableResult <= {9'b010111111};
9'b001000000: tableResult <= {9'b100000000};
9'b001000001: tableResult <= {9'b100000100};
9'b001000010: tableResult <= {9'b010000100};
9'b001000011: tableResult <= {9'b001000100};
9'b001000100: tableResult <= {9'b001000100};
9'b001000101: tableResult <= {9'b000000100};
9'b001000110: tableResult <= {9'b010010111};
9'b001000111: tableResult <= {9'b010010111};
9'b001001000: tableResult <= {9'b100100000};
9'b001001001: tableResult <= {9'b010010010};
9'b001001010: tableResult <= {9'b001001010};
9'b001001011: tableResult <= {9'b001001011};
9'b001001100: tableResult <= {9'b001001011};
9'b001001101: tableResult <= {9'b010011111};
9'b001001110: tableResult <= {9'b010011111};
9'b001001111: tableResult <= {9'b010011111};
9'b001010000: tableResult <= {9'b010100000};
9'b001010001: tableResult <= {9'b001010001};
9'b001010010: tableResult <= {9'b001010010};
9'b001010011: tableResult <= {9'b001010011};
9'b001010100: tableResult <= {9'b001001011};
9'b001010101: tableResult <= {9'b010011111};
9'b001010110: tableResult <= {9'b010011111};
9'b001010111: tableResult <= {9'b010011111};
9'b001011000: tableResult <= {9'b001100000};
9'b001011001: tableResult <= {9'b001011001};
9'b001011010: tableResult <= {9'b001011010};
9'b001011011: tableResult <= {9'b001011011};
9'b001011100: tableResult <= {9'b001010011};
9'b001011101: tableResult <= {9'b010100111};
9'b001011110: tableResult <= {9'b010100111};
9'b001011111: tableResult <= {9'b010011111};
9'b001100000: tableResult <= {9'b001100000};
9'b001100001: tableResult <= {9'b001011001};
9'b001100010: tableResult <= {9'b001011001};
9'b001100011: tableResult <= {9'b001011010};
9'b001100100: tableResult <= {9'b001011011};
9'b001100101: tableResult <= {9'b010110111};
9'b001100110: tableResult <= {9'b010101111};
9'b001100111: tableResult <= {9'b010100111};
9'b001101000: tableResult <= {9'b000100000};
9'b001101001: tableResult <= {9'b010111011};
9'b001101010: tableResult <= {9'b010111011};
9'b001101011: tableResult <= {9'b010111100};
9'b001101100: tableResult <= {9'b010111110};
9'b001101101: tableResult <= {9'b010111111};
9'b001101110: tableResult <= {9'b010110111};
9'b001101111: tableResult <= {9'b010101111};
9'b001110000: tableResult <= {9'b010111010};
9'b001110001: tableResult <= {9'b010111011};
9'b001110010: tableResult <= {9'b010111011};
9'b001110011: tableResult <= {9'b010111100};
9'b001110100: tableResult <= {9'b010111101};
9'b001110101: tableResult <= {9'b010111110};
9'b001110110: tableResult <= {9'b010111111};
9'b001110111: tableResult <= {9'b010110111};
9'b001111000: tableResult <= {9'b010111010};
9'b001111001: tableResult <= {9'b010111011};
9'b001111010: tableResult <= {9'b010111011};
9'b001111011: tableResult <= {9'b010111011};
9'b001111100: tableResult <= {9'b010111100};
9'b001111101: tableResult <= {9'b010111101};
9'b001111110: tableResult <= {9'b010111110};
9'b001111111: tableResult <= {9'b010111111};
9'b010000000: tableResult <= {9'b100000000};
9'b010000001: tableResult <= {9'b100000010};
9'b010000010: tableResult <= {9'b100000100};
9'b010000011: tableResult <= {9'b011000100};
9'b010000100: tableResult <= {9'b010000100};
9'b010000101: tableResult <= {9'b001000100};
9'b010000110: tableResult <= {9'b011010111};
9'b010000111: tableResult <= {9'b011010111};
9'b010001000: tableResult <= {9'b100010000};
9'b010001001: tableResult <= {9'b010001001};
9'b010001010: tableResult <= {9'b010001010};
9'b010001011: tableResult <= {9'b010001011};
9'b010001100: tableResult <= {9'b001001011};
9'b010001101: tableResult <= {9'b100010111};
9'b010001110: tableResult <= {9'b011010111};
9'b010001111: tableResult <= {9'b011010111};
9'b010010000: tableResult <= {9'b100100000};
9'b010010001: tableResult <= {9'b010010001};
9'b010010010: tableResult <= {9'b010010010};
9'b010010011: tableResult <= {9'b001001010};
9'b010010100: tableResult <= {9'b100100101};
9'b010010101: tableResult <= {9'b011011110};
9'b010010110: tableResult <= {9'b011011110};
9'b010010111: tableResult <= {9'b010011111};
9'b010011000: tableResult <= {9'b011100000};
9'b010011001: tableResult <= {9'b010011001};
9'b010011010: tableResult <= {9'b001010001};
9'b010011011: tableResult <= {9'b001010010};
9'b010011100: tableResult <= {9'b100100101};
9'b010011101: tableResult <= {9'b011100110};
9'b010011110: tableResult <= {9'b011100110};
9'b010011111: tableResult <= {9'b010011111};
9'b010100000: tableResult <= {9'b010100000};
9'b010100001: tableResult <= {9'b001011001};
9'b010100010: tableResult <= {9'b100101100};
9'b010100011: tableResult <= {9'b100101100};
9'b010100100: tableResult <= {9'b100101101};
9'b010100101: tableResult <= {9'b011101110};
9'b010100110: tableResult <= {9'b011100110};
9'b010100111: tableResult <= {9'b010100111};
9'b010101000: tableResult <= {9'b001100000};
9'b010101001: tableResult <= {9'b100111010};
9'b010101010: tableResult <= {9'b011110011};
9'b010101011: tableResult <= {9'b011110100};
9'b010101100: tableResult <= {9'b011110101};
9'b010101101: tableResult <= {9'b011110110};
9'b010101110: tableResult <= {9'b011101110};
9'b010101111: tableResult <= {9'b010101111};
9'b010110000: tableResult <= {9'b011111010};
9'b010110001: tableResult <= {9'b011111010};
9'b010110010: tableResult <= {9'b011110011};
9'b010110011: tableResult <= {9'b011110100};
9'b010110100: tableResult <= {9'b011110100};
9'b010110101: tableResult <= {9'b011110101};
9'b010110110: tableResult <= {9'b011110110};
9'b010110111: tableResult <= {9'b010110111};
9'b010111000: tableResult <= {9'b011111010};
9'b010111001: tableResult <= {9'b011111010};
9'b010111010: tableResult <= {9'b010111011};
9'b010111011: tableResult <= {9'b010111011};
9'b010111100: tableResult <= {9'b010111100};
9'b010111101: tableResult <= {9'b010111101};
9'b010111110: tableResult <= {9'b010111110};
9'b010111111: tableResult <= {9'b010111111};
9'b011000000: tableResult <= {9'b100000000};
9'b011000001: tableResult <= {9'b100000001};
9'b011000010: tableResult <= {9'b100000011};
9'b011000011: tableResult <= {9'b100000100};
9'b011000100: tableResult <= {9'b011000100};
9'b011000101: tableResult <= {9'b011000100};
9'b011000110: tableResult <= {9'b101010111};
9'b011000111: tableResult <= {9'b101010111};
9'b011001000: tableResult <= {9'b100001000};
9'b011001001: tableResult <= {9'b011001001};
9'b011001010: tableResult <= {9'b011001010};
9'b011001011: tableResult <= {9'b011001011};
9'b011001100: tableResult <= {9'b010001011};
9'b011001101: tableResult <= {9'b101010111};
9'b011001110: tableResult <= {9'b100010111};
9'b011001111: tableResult <= {9'b100010111};
9'b011010000: tableResult <= {9'b100011000};
9'b011010001: tableResult <= {9'b011010001};
9'b011010010: tableResult <= {9'b010001001};
9'b011010011: tableResult <= {9'b010001010};
9'b011010100: tableResult <= {9'b101100101};
9'b011010101: tableResult <= {9'b100011110};
9'b011010110: tableResult <= {9'b100011110};
9'b011010111: tableResult <= {9'b011010111};
9'b011011000: tableResult <= {9'b100100000};
9'b011011001: tableResult <= {9'b011011001};
9'b011011010: tableResult <= {9'b010010001};
9'b011011011: tableResult <= {9'b101101101};
9'b011011100: tableResult <= {9'b100100101};
9'b011011101: tableResult <= {9'b100100101};
9'b011011110: tableResult <= {9'b011011110};
9'b011011111: tableResult <= {9'b010011111};
9'b011100000: tableResult <= {9'b011100000};
9'b011100001: tableResult <= {9'b010011001};
9'b011100010: tableResult <= {9'b101101100};
9'b011100011: tableResult <= {9'b100101100};
9'b011100100: tableResult <= {9'b100101101};
9'b011100101: tableResult <= {9'b100100101};
9'b011100110: tableResult <= {9'b011100110};
9'b011100111: tableResult <= {9'b010011111};
9'b011101000: tableResult <= {9'b011100000};
9'b011101001: tableResult <= {9'b101111010};
9'b011101010: tableResult <= {9'b100110011};
9'b011101011: tableResult <= {9'b100101100};
9'b011101100: tableResult <= {9'b100101100};
9'b011101101: tableResult <= {9'b100101101};
9'b011101110: tableResult <= {9'b011101110};
9'b011101111: tableResult <= {9'b010100111};
9'b011110000: tableResult <= {9'b101111010};
9'b011110001: tableResult <= {9'b100111010};
9'b011110010: tableResult <= {9'b100110011};
9'b011110011: tableResult <= {9'b011110011};
9'b011110100: tableResult <= {9'b011110100};
9'b011110101: tableResult <= {9'b011110101};
9'b011110110: tableResult <= {9'b011110110};
9'b011110111: tableResult <= {9'b010110111};
9'b011111000: tableResult <= {9'b101111010};
9'b011111001: tableResult <= {9'b100111010};
9'b011111010: tableResult <= {9'b011111010};
9'b011111011: tableResult <= {9'b010111011};
9'b011111100: tableResult <= {9'b010111011};
9'b011111101: tableResult <= {9'b010111100};
9'b011111110: tableResult <= {9'b010111110};
9'b011111111: tableResult <= {9'b010111111};
9'b100000000: tableResult <= {9'b100000000};
9'b100000001: tableResult <= {9'b100000000};
9'b100000010: tableResult <= {9'b100000010};
9'b100000011: tableResult <= {9'b100000011};
9'b100000100: tableResult <= {9'b100000100};
9'b100000101: tableResult <= {9'b100000100};
9'b100000110: tableResult <= {9'b110010111};
9'b100000111: tableResult <= {9'b101010111};
9'b100001000: tableResult <= {9'b100000000};
9'b100001001: tableResult <= {9'b011001001};
9'b100001010: tableResult <= {9'b011001010};
9'b100001011: tableResult <= {9'b011001010};
9'b100001100: tableResult <= {9'b011001011};
9'b100001101: tableResult <= {9'b101010111};
9'b100001110: tableResult <= {9'b101010111};
9'b100001111: tableResult <= {9'b101010111};
9'b100010000: tableResult <= {9'b100010000};
9'b100010001: tableResult <= {9'b011010001};
9'b100010010: tableResult <= {9'b101100100};
9'b100010011: tableResult <= {9'b101100101};
9'b100010100: tableResult <= {9'b101100101};
9'b100010101: tableResult <= {9'b101011110};
9'b100010110: tableResult <= {9'b101011110};
9'b100010111: tableResult <= {9'b100010111};
9'b100011000: tableResult <= {9'b100011000};
9'b100011001: tableResult <= {9'b011010001};
9'b100011010: tableResult <= {9'b101101100};
9'b100011011: tableResult <= {9'b101100100};
9'b100011100: tableResult <= {9'b101100101};
9'b100011101: tableResult <= {9'b101100101};
9'b100011110: tableResult <= {9'b100011110};
9'b100011111: tableResult <= {9'b100010111};
9'b100100000: tableResult <= {9'b100100000};
9'b100100001: tableResult <= {9'b011011001};
9'b100100010: tableResult <= {9'b101101100};
9'b100100011: tableResult <= {9'b101101100};
9'b100100100: tableResult <= {9'b101101101};
9'b100100101: tableResult <= {9'b100100101};
9'b100100110: tableResult <= {9'b100100101};
9'b100100111: tableResult <= {9'b111111111};
9'b100101000: tableResult <= {9'b100100000};
9'b100101001: tableResult <= {9'b101111010};
9'b100101010: tableResult <= {9'b101110011};
9'b100101011: tableResult <= {9'b101101100};
9'b100101100: tableResult <= {9'b100101100};
9'b100101101: tableResult <= {9'b100101101};
9'b100101110: tableResult <= {9'b100100101};
9'b100101111: tableResult <= {9'b111111111};
9'b100110000: tableResult <= {9'b110111010};
9'b100110001: tableResult <= {9'b101111010};
9'b100110010: tableResult <= {9'b101110011};
9'b100110011: tableResult <= {9'b100110011};
9'b100110100: tableResult <= {9'b100101100};
9'b100110101: tableResult <= {9'b100101100};
9'b100110110: tableResult <= {9'b100101101};
9'b100110111: tableResult <= {9'b111111111};
9'b100111000: tableResult <= {9'b101111010};
9'b100111001: tableResult <= {9'b101111010};
9'b100111010: tableResult <= {9'b100111010};
9'b100111011: tableResult <= {9'b100111010};
9'b100111100: tableResult <= {9'b111111111};
9'b100111101: tableResult <= {9'b111111111};
9'b100111110: tableResult <= {9'b111111111};
9'b100111111: tableResult <= {9'b111111111};
9'b101000000: tableResult <= {9'b100000000};
9'b101000001: tableResult <= {9'b100000000};
9'b101000010: tableResult <= {9'b100000001};
9'b101000011: tableResult <= {9'b100000010};
9'b101000100: tableResult <= {9'b100000011};
9'b101000101: tableResult <= {9'b100000100};
9'b101000110: tableResult <= {9'b111010111};
9'b101000111: tableResult <= {9'b110010111};
9'b101001000: tableResult <= {9'b100000000};
9'b101001001: tableResult <= {9'b111010010};
9'b101001010: tableResult <= {9'b111010011};
9'b101001011: tableResult <= {9'b111010101};
9'b101001100: tableResult <= {9'b111010110};
9'b101001101: tableResult <= {9'b111010110};
9'b101001110: tableResult <= {9'b110010111};
9'b101001111: tableResult <= {9'b101010111};
9'b101010000: tableResult <= {9'b100001000};
9'b101010001: tableResult <= {9'b111011010};
9'b101010010: tableResult <= {9'b110011011};
9'b101010011: tableResult <= {9'b110011100};
9'b101010100: tableResult <= {9'b110011101};
9'b101010101: tableResult <= {9'b110011110};
9'b101010110: tableResult <= {9'b101011110};
9'b101010111: tableResult <= {9'b101010111};
9'b101011000: tableResult <= {9'b100010000};
9'b101011001: tableResult <= {9'b111101010};
9'b101011010: tableResult <= {9'b110100011};
9'b101011011: tableResult <= {9'b101100100};
9'b101011100: tableResult <= {9'b101100101};
9'b101011101: tableResult <= {9'b101100101};
9'b101011110: tableResult <= {9'b101011110};
9'b101011111: tableResult <= {9'b101010111};
9'b101100000: tableResult <= {9'b100011000};
9'b101100001: tableResult <= {9'b111110010};
9'b101100010: tableResult <= {9'b110101011};
9'b101100011: tableResult <= {9'b101101100};
9'b101100100: tableResult <= {9'b101100100};
9'b101100101: tableResult <= {9'b101100101};
9'b101100110: tableResult <= {9'b101100101};
9'b101100111: tableResult <= {9'b111111111};
9'b101101000: tableResult <= {9'b100100000};
9'b101101001: tableResult <= {9'b111110010};
9'b101101010: tableResult <= {9'b110110011};
9'b101101011: tableResult <= {9'b101101100};
9'b101101100: tableResult <= {9'b101101100};
9'b101101101: tableResult <= {9'b101101101};
9'b101101110: tableResult <= {9'b111111111};
9'b101101111: tableResult <= {9'b111111111};
9'b101110000: tableResult <= {9'b111111010};
9'b101110001: tableResult <= {9'b110111010};
9'b101110010: tableResult <= {9'b101110011};
9'b101110011: tableResult <= {9'b101110011};
9'b101110100: tableResult <= {9'b101101100};
9'b101110101: tableResult <= {9'b111111111};
9'b101110110: tableResult <= {9'b111111111};
9'b101110111: tableResult <= {9'b111111111};
9'b101111000: tableResult <= {9'b110111010};
9'b101111001: tableResult <= {9'b101111010};
9'b101111010: tableResult <= {9'b101111010};
9'b101111011: tableResult <= {9'b101111010};
9'b101111100: tableResult <= {9'b111111111};
9'b101111101: tableResult <= {9'b111111111};
9'b101111110: tableResult <= {9'b111111111};
9'b101111111: tableResult <= {9'b111111111};
9'b110000000: tableResult <= {9'b111010010};
9'b110000001: tableResult <= {9'b111010011};
9'b110000010: tableResult <= {9'b111010100};
9'b110000011: tableResult <= {9'b111010101};
9'b110000100: tableResult <= {9'b111010110};
9'b110000101: tableResult <= {9'b111010110};
9'b110000110: tableResult <= {9'b111010111};
9'b110000111: tableResult <= {9'b111010111};
9'b110001000: tableResult <= {9'b111011010};
9'b110001001: tableResult <= {9'b111010010};
9'b110001010: tableResult <= {9'b111010011};
9'b110001011: tableResult <= {9'b111010100};
9'b110001100: tableResult <= {9'b111010101};
9'b110001101: tableResult <= {9'b111010110};
9'b110001110: tableResult <= {9'b111010110};
9'b110001111: tableResult <= {9'b110010111};
9'b110010000: tableResult <= {9'b111100010};
9'b110010001: tableResult <= {9'b111011010};
9'b110010010: tableResult <= {9'b110011011};
9'b110010011: tableResult <= {9'b110011100};
9'b110010100: tableResult <= {9'b110011101};
9'b110010101: tableResult <= {9'b110011101};
9'b110010110: tableResult <= {9'b110011110};
9'b110010111: tableResult <= {9'b110010111};
9'b110011000: tableResult <= {9'b111101010};
9'b110011001: tableResult <= {9'b111100010};
9'b110011010: tableResult <= {9'b110100011};
9'b110011011: tableResult <= {9'b110011011};
9'b110011100: tableResult <= {9'b110011100};
9'b110011101: tableResult <= {9'b110011101};
9'b110011110: tableResult <= {9'b110011110};
9'b110011111: tableResult <= {9'b101010111};
9'b110100000: tableResult <= {9'b111110010};
9'b110100001: tableResult <= {9'b111101010};
9'b110100010: tableResult <= {9'b110101011};
9'b110100011: tableResult <= {9'b110100011};
9'b110100100: tableResult <= {9'b101100100};
9'b110100101: tableResult <= {9'b101100101};
9'b110100110: tableResult <= {9'b101100101};
9'b110100111: tableResult <= {9'b111111111};
9'b110101000: tableResult <= {9'b111110010};
9'b110101001: tableResult <= {9'b111110010};
9'b110101010: tableResult <= {9'b110101011};
9'b110101011: tableResult <= {9'b110101011};
9'b110101100: tableResult <= {9'b101101100};
9'b110101101: tableResult <= {9'b111111111};
9'b110101110: tableResult <= {9'b111111111};
9'b110101111: tableResult <= {9'b111111111};
9'b110110000: tableResult <= {9'b111111010};
9'b110110001: tableResult <= {9'b111110010};
9'b110110010: tableResult <= {9'b110110011};
9'b110110011: tableResult <= {9'b110110011};
9'b110110100: tableResult <= {9'b101101100};
9'b110110101: tableResult <= {9'b111111111};
9'b110110110: tableResult <= {9'b111111111};
9'b110110111: tableResult <= {9'b111111111};
9'b110111000: tableResult <= {9'b111111010};
9'b110111001: tableResult <= {9'b110111010};
9'b110111010: tableResult <= {9'b110111010};
9'b110111011: tableResult <= {9'b101111010};
9'b110111100: tableResult <= {9'b111111111};
9'b110111101: tableResult <= {9'b111111111};
9'b110111110: tableResult <= {9'b111111111};
9'b110111111: tableResult <= {9'b111111111};
9'b111000000: tableResult <= {9'b111010010};
9'b111000001: tableResult <= {9'b111010011};
9'b111000010: tableResult <= {9'b111010100};
9'b111000011: tableResult <= {9'b111010100};
9'b111000100: tableResult <= {9'b111010101};
9'b111000101: tableResult <= {9'b111010110};
9'b111000110: tableResult <= {9'b111010111};
9'b111000111: tableResult <= {9'b111010111};
9'b111001000: tableResult <= {9'b111011010};
9'b111001001: tableResult <= {9'b111010010};
9'b111001010: tableResult <= {9'b111010011};
9'b111001011: tableResult <= {9'b111010100};
9'b111001100: tableResult <= {9'b111010101};
9'b111001101: tableResult <= {9'b111010110};
9'b111001110: tableResult <= {9'b111010110};
9'b111001111: tableResult <= {9'b111010110};
9'b111010000: tableResult <= {9'b111100010};
9'b111010001: tableResult <= {9'b111011010};
9'b111010010: tableResult <= {9'b111010010};
9'b111010011: tableResult <= {9'b111010011};
9'b111010100: tableResult <= {9'b111010100};
9'b111010101: tableResult <= {9'b111010101};
9'b111010110: tableResult <= {9'b111010110};
9'b111010111: tableResult <= {9'b111010110};
9'b111011000: tableResult <= {9'b111100010};
9'b111011001: tableResult <= {9'b111100010};
9'b111011010: tableResult <= {9'b111011010};
9'b111011011: tableResult <= {9'b111010010};
9'b111011100: tableResult <= {9'b111010011};
9'b111011101: tableResult <= {9'b111010101};
9'b111011110: tableResult <= {9'b111010110};
9'b111011111: tableResult <= {9'b111010110};
9'b111100000: tableResult <= {9'b111101010};
9'b111100001: tableResult <= {9'b111101010};
9'b111100010: tableResult <= {9'b111100010};
9'b111100011: tableResult <= {9'b111011010};
9'b111100100: tableResult <= {9'b111111111};
9'b111100101: tableResult <= {9'b111111111};
9'b111100110: tableResult <= {9'b111111111};
9'b111100111: tableResult <= {9'b111111111};
9'b111101000: tableResult <= {9'b111110010};
9'b111101001: tableResult <= {9'b111110010};
9'b111101010: tableResult <= {9'b111101010};
9'b111101011: tableResult <= {9'b111101010};
9'b111101100: tableResult <= {9'b111111111};
9'b111101101: tableResult <= {9'b111111111};
9'b111101110: tableResult <= {9'b111111111};
9'b111101111: tableResult <= {9'b111111111};
9'b111110000: tableResult <= {9'b111111010};
9'b111110001: tableResult <= {9'b111110010};
9'b111110010: tableResult <= {9'b111110010};
9'b111110011: tableResult <= {9'b111110010};
9'b111110100: tableResult <= {9'b111111111};
9'b111110101: tableResult <= {9'b111111111};
9'b111110110: tableResult <= {9'b111111111};
9'b111110111: tableResult <= {9'b111111111};
9'b111111000: tableResult <= {9'b111111010};
9'b111111001: tableResult <= {9'b111110010};
9'b111111010: tableResult <= {9'b111110010};
9'b111111011: tableResult <= {9'b111110010};
9'b111111100: tableResult <= {9'b111111111};
9'b111111101: tableResult <= {9'b111111111};
9'b111111110: tableResult <= {9'b111111111};
9'b111111111: tableResult <= {9'b111111111};
			//end code from matlab
			default: tableResult <= 9'd0;
		endcase
	end
	
endmodule
