/****************************************************************
 * Skyler Schneider ss868                                       *
 * ECE 5760 Final Project                                       *
 * Sand Game                                                    *
 ****************************************************************/

// ROM that stores the pixel data for the troll images. Each word
// of 16 bits stores eight 2-bit pixel data. There are four pictures
// in the animation, each 160 pixels wide by 120 pixels high.
module TrollROM (
    input             iCLK,  // Clock signal for reading
    input      [13:0] iAddr, // (Pic# * 2400) + (Y * 20) + (X/8)
    output reg [15:0] oData  // Pixel value (actually 8 pixels)
);
    
    always @(posedge iCLK) begin
        case(iAddr)
            14'h0000: oData <= 16'h0000;
            14'h0001: oData <= 16'h0000;
            14'h0002: oData <= 16'h0000;
            14'h0003: oData <= 16'ha800;
            14'h0004: oData <= 16'h0000;
            14'h0005: oData <= 16'h0000;
            14'h0006: oData <= 16'h0000;
            14'h0007: oData <= 16'h0000;
            14'h0008: oData <= 16'h0000;
            14'h0009: oData <= 16'h0000;
            14'h000a: oData <= 16'h0000;
            14'h000b: oData <= 16'h0000;
            14'h000c: oData <= 16'h0000;
            14'h000d: oData <= 16'h0000;
            14'h000e: oData <= 16'h0000;
            14'h000f: oData <= 16'h0000;
            14'h0010: oData <= 16'h0000;
            14'h0011: oData <= 16'h0000;
            14'h0012: oData <= 16'h0000;
            14'h0013: oData <= 16'h0000;
            14'h0014: oData <= 16'h0000;
            14'h0015: oData <= 16'h0000;
            14'h0016: oData <= 16'h0000;
            14'h0017: oData <= 16'haa00;
            14'h0018: oData <= 16'h0002;
            14'h0019: oData <= 16'h0000;
            14'h001a: oData <= 16'ha800;
            14'h001b: oData <= 16'haaaa;
            14'h001c: oData <= 16'haaaa;
            14'h001d: oData <= 16'haaaa;
            14'h001e: oData <= 16'haaaa;
            14'h001f: oData <= 16'h0002;
            14'h0020: oData <= 16'h0000;
            14'h0021: oData <= 16'h0000;
            14'h0022: oData <= 16'h0000;
            14'h0023: oData <= 16'h0000;
            14'h0024: oData <= 16'h0000;
            14'h0025: oData <= 16'h0000;
            14'h0026: oData <= 16'h0000;
            14'h0027: oData <= 16'h0000;
            14'h0028: oData <= 16'h0000;
            14'h0029: oData <= 16'h0000;
            14'h002a: oData <= 16'h0000;
            14'h002b: oData <= 16'haa00;
            14'h002c: oData <= 16'h0002;
            14'h002d: oData <= 16'h0000;
            14'h002e: oData <= 16'haa80;
            14'h002f: oData <= 16'haaaa;
            14'h0030: oData <= 16'haaaa;
            14'h0031: oData <= 16'haaaa;
            14'h0032: oData <= 16'haaaa;
            14'h0033: oData <= 16'haaaa;
            14'h0034: oData <= 16'h00aa;
            14'h0035: oData <= 16'h0000;
            14'h0036: oData <= 16'h0000;
            14'h0037: oData <= 16'h0000;
            14'h0038: oData <= 16'h0000;
            14'h0039: oData <= 16'h0000;
            14'h003a: oData <= 16'h0000;
            14'h003b: oData <= 16'h0000;
            14'h003c: oData <= 16'h0000;
            14'h003d: oData <= 16'h0000;
            14'h003e: oData <= 16'h0000;
            14'h003f: oData <= 16'ha800;
            14'h0040: oData <= 16'h000a;
            14'h0041: oData <= 16'h0000;
            14'h0042: oData <= 16'hfaa8;
            14'h0043: oData <= 16'hffff;
            14'h0044: oData <= 16'hffff;
            14'h0045: oData <= 16'hffff;
            14'h0046: oData <= 16'hffff;
            14'h0047: oData <= 16'haaaa;
            14'h0048: oData <= 16'haaaa;
            14'h0049: oData <= 16'h0000;
            14'h004a: oData <= 16'h0000;
            14'h004b: oData <= 16'h0000;
            14'h004c: oData <= 16'h0000;
            14'h004d: oData <= 16'h0000;
            14'h004e: oData <= 16'h0000;
            14'h004f: oData <= 16'h0000;
            14'h0050: oData <= 16'h0000;
            14'h0051: oData <= 16'h0000;
            14'h0052: oData <= 16'h0aa8;
            14'h0053: oData <= 16'ha800;
            14'h0054: oData <= 16'h000a;
            14'h0055: oData <= 16'h0000;
            14'h0056: oData <= 16'hffaa;
            14'h0057: oData <= 16'hffff;
            14'h0058: oData <= 16'haabf;
            14'h0059: oData <= 16'haaaa;
            14'h005a: oData <= 16'hffaa;
            14'h005b: oData <= 16'hffff;
            14'h005c: oData <= 16'haabf;
            14'h005d: oData <= 16'h02aa;
            14'h005e: oData <= 16'h0000;
            14'h005f: oData <= 16'h0000;
            14'h0060: oData <= 16'h0000;
            14'h0061: oData <= 16'h0000;
            14'h0062: oData <= 16'h0000;
            14'h0063: oData <= 16'h0000;
            14'h0064: oData <= 16'h0000;
            14'h0065: oData <= 16'h0000;
            14'h0066: oData <= 16'haaaa;
            14'h0067: oData <= 16'ha002;
            14'h0068: oData <= 16'h002a;
            14'h0069: oData <= 16'h8000;
            14'h006a: oData <= 16'hfffa;
            14'h006b: oData <= 16'hffff;
            14'h006c: oData <= 16'hffea;
            14'h006d: oData <= 16'hffff;
            14'h006e: oData <= 16'haaff;
            14'h006f: oData <= 16'haaaa;
            14'h0070: oData <= 16'hbfaa;
            14'h0071: oData <= 16'h2aaa;
            14'h0072: oData <= 16'h0000;
            14'h0073: oData <= 16'h0000;
            14'h0074: oData <= 16'h0000;
            14'h0075: oData <= 16'h0000;
            14'h0076: oData <= 16'h0000;
            14'h0077: oData <= 16'h0000;
            14'h0078: oData <= 16'h0000;
            14'h0079: oData <= 16'h0000;
            14'h007a: oData <= 16'haaaa;
            14'h007b: oData <= 16'ha00a;
            14'h007c: oData <= 16'h002a;
            14'h007d: oData <= 16'ha00a;
            14'h007e: oData <= 16'hfffe;
            14'h007f: oData <= 16'hafff;
            14'h0080: oData <= 16'hffff;
            14'h0081: oData <= 16'heaaa;
            14'h0082: oData <= 16'hffff;
            14'h0083: oData <= 16'hffff;
            14'h0084: oData <= 16'hffff;
            14'h0085: oData <= 16'haaff;
            14'h0086: oData <= 16'h0000;
            14'h0087: oData <= 16'h0000;
            14'h0088: oData <= 16'h0000;
            14'h0089: oData <= 16'h0000;
            14'h008a: oData <= 16'h0000;
            14'h008b: oData <= 16'h0000;
            14'h008c: oData <= 16'h0000;
            14'h008d: oData <= 16'h8000;
            14'h008e: oData <= 16'haaaa;
            14'h008f: oData <= 16'h802a;
            14'h0090: oData <= 16'ha0aa;
            14'h0091: oData <= 16'ha02a;
            14'h0092: oData <= 16'hffff;
            14'h0093: oData <= 16'hfaff;
            14'h0094: oData <= 16'haabf;
            14'h0095: oData <= 16'hbfff;
            14'h0096: oData <= 16'hffea;
            14'h0097: oData <= 16'hffff;
            14'h0098: oData <= 16'haaff;
            14'h0099: oData <= 16'haffa;
            14'h009a: oData <= 16'h000a;
            14'h009b: oData <= 16'h0000;
            14'h009c: oData <= 16'h0000;
            14'h009d: oData <= 16'h0000;
            14'h009e: oData <= 16'h0000;
            14'h009f: oData <= 16'h0000;
            14'h00a0: oData <= 16'h0000;
            14'h00a1: oData <= 16'ha000;
            14'h00a2: oData <= 16'haaaa;
            14'h00a3: oData <= 16'h80aa;
            14'h00a4: oData <= 16'ha8aa;
            14'h00a5: oData <= 16'ha82a;
            14'h00a6: oData <= 16'hffff;
            14'h00a7: oData <= 16'hffaf;
            14'h00a8: oData <= 16'hffea;
            14'h00a9: oData <= 16'hffff;
            14'h00aa: oData <= 16'haabf;
            14'h00ab: oData <= 16'haaaa;
            14'h00ac: oData <= 16'hffaa;
            14'h00ad: oData <= 16'hbfaf;
            14'h00ae: oData <= 16'h00aa;
            14'h00af: oData <= 16'h0000;
            14'h00b0: oData <= 16'h0000;
            14'h00b1: oData <= 16'h0000;
            14'h00b2: oData <= 16'h0000;
            14'h00b3: oData <= 16'h0000;
            14'h00b4: oData <= 16'h0000;
            14'h00b5: oData <= 16'ha000;
            14'h00b6: oData <= 16'h802a;
            14'h00b7: oData <= 16'h00aa;
            14'h00b8: oData <= 16'haaaa;
            14'h00b9: oData <= 16'hea2a;
            14'h00ba: oData <= 16'hffff;
            14'h00bb: oData <= 16'haffa;
            14'h00bc: oData <= 16'hafff;
            14'h00bd: oData <= 16'haaaa;
            14'h00be: oData <= 16'hffff;
            14'h00bf: oData <= 16'hffff;
            14'h00c0: oData <= 16'hffff;
            14'h00c1: oData <= 16'hffbf;
            14'h00c2: oData <= 16'h02ab;
            14'h00c3: oData <= 16'h0000;
            14'h00c4: oData <= 16'h0000;
            14'h00c5: oData <= 16'h0000;
            14'h00c6: oData <= 16'h0000;
            14'h00c7: oData <= 16'h0000;
            14'h00c8: oData <= 16'h0000;
            14'h00c9: oData <= 16'ha000;
            14'h00ca: oData <= 16'h000a;
            14'h00cb: oData <= 16'h02aa;
            14'h00cc: oData <= 16'haaaa;
            14'h00cd: oData <= 16'hfa8a;
            14'h00ce: oData <= 16'hbfff;
            14'h00cf: oData <= 16'hfaff;
            14'h00d0: oData <= 16'hfaaf;
            14'h00d1: oData <= 16'hbfff;
            14'h00d2: oData <= 16'hfffe;
            14'h00d3: oData <= 16'hffff;
            14'h00d4: oData <= 16'haabf;
            14'h00d5: oData <= 16'hffff;
            14'h00d6: oData <= 16'h0abf;
            14'h00d7: oData <= 16'h0000;
            14'h00d8: oData <= 16'h0000;
            14'h00d9: oData <= 16'h0000;
            14'h00da: oData <= 16'h0000;
            14'h00db: oData <= 16'h0000;
            14'h00dc: oData <= 16'h0000;
            14'h00dd: oData <= 16'ha800;
            14'h00de: oData <= 16'h000a;
            14'h00df: oData <= 16'h02aa;
            14'h00e0: oData <= 16'haaa8;
            14'h00e1: oData <= 16'hfe80;
            14'h00e2: oData <= 16'hebff;
            14'h00e3: oData <= 16'hbfaf;
            14'h00e4: oData <= 16'hfffa;
            14'h00e5: oData <= 16'hebff;
            14'h00e6: oData <= 16'hffff;
            14'h00e7: oData <= 16'hafff;
            14'h00e8: oData <= 16'hbfea;
            14'h00e9: oData <= 16'hfffe;
            14'h00ea: oData <= 16'h2aff;
            14'h00eb: oData <= 16'h0000;
            14'h00ec: oData <= 16'h0000;
            14'h00ed: oData <= 16'h0000;
            14'h00ee: oData <= 16'h0000;
            14'h00ef: oData <= 16'h0000;
            14'h00f0: oData <= 16'h0000;
            14'h00f1: oData <= 16'ha800;
            14'h00f2: oData <= 16'h000a;
            14'h00f3: oData <= 16'h02a8;
            14'h00f4: oData <= 16'h2aa0;
            14'h00f5: oData <= 16'hfea0;
            14'h00f6: oData <= 16'hfeff;
            14'h00f7: oData <= 16'hebfb;
            14'h00f8: oData <= 16'hffff;
            14'h00f9: oData <= 16'hafff;
            14'h00fa: oData <= 16'hffff;
            14'h00fb: oData <= 16'hfabf;
            14'h00fc: oData <= 16'hffff;
            14'h00fd: oData <= 16'hffeb;
            14'h00fe: oData <= 16'h2bff;
            14'h00ff: oData <= 16'h0000;
            14'h0100: oData <= 16'h0000;
            14'h0101: oData <= 16'h0000;
            14'h0102: oData <= 16'h0000;
            14'h0103: oData <= 16'h0000;
            14'h0104: oData <= 16'h0000;
            14'h0105: oData <= 16'ha800;
            14'h0106: oData <= 16'h000a;
            14'h0107: oData <= 16'h02a8;
            14'h0108: oData <= 16'h2aa0;
            14'h0109: oData <= 16'hffa0;
            14'h010a: oData <= 16'hffbf;
            14'h010b: oData <= 16'hfefe;
            14'h010c: oData <= 16'hffff;
            14'h010d: oData <= 16'hbfff;
            14'h010e: oData <= 16'hffff;
            14'h010f: oData <= 16'hffbf;
            14'h0110: oData <= 16'hffff;
            14'h0111: oData <= 16'hffbf;
            14'h0112: oData <= 16'h2bff;
            14'h0113: oData <= 16'h0000;
            14'h0114: oData <= 16'h0000;
            14'h0115: oData <= 16'h0000;
            14'h0116: oData <= 16'h0000;
            14'h0117: oData <= 16'h0000;
            14'h0118: oData <= 16'h00a8;
            14'h0119: oData <= 16'ha800;
            14'h011a: oData <= 16'h000a;
            14'h011b: oData <= 16'h02a8;
            14'h011c: oData <= 16'h0a80;
            14'h011d: oData <= 16'hffa0;
            14'h011e: oData <= 16'hbfff;
            14'h011f: oData <= 16'hffbf;
            14'h0120: oData <= 16'hffff;
            14'h0121: oData <= 16'hbfff;
            14'h0122: oData <= 16'hfffe;
            14'h0123: oData <= 16'hefff;
            14'h0124: oData <= 16'hffff;
            14'h0125: oData <= 16'hffbf;
            14'h0126: oData <= 16'h2bff;
            14'h0127: oData <= 16'h0000;
            14'h0128: oData <= 16'h0000;
            14'h0129: oData <= 16'h0000;
            14'h012a: oData <= 16'h0000;
            14'h012b: oData <= 16'h0000;
            14'h012c: oData <= 16'h02aa;
            14'h012d: oData <= 16'ha000;
            14'h012e: oData <= 16'h000a;
            14'h012f: oData <= 16'h02a8;
            14'h0130: oData <= 16'h0000;
            14'h0131: oData <= 16'hffa8;
            14'h0132: oData <= 16'hefff;
            14'h0133: oData <= 16'hffef;
            14'h0134: oData <= 16'hffff;
            14'h0135: oData <= 16'hffff;
            14'h0136: oData <= 16'hfffe;
            14'h0137: oData <= 16'hfbff;
            14'h0138: oData <= 16'hffff;
            14'h0139: oData <= 16'hfeff;
            14'h013a: oData <= 16'h2bff;
            14'h013b: oData <= 16'h0000;
            14'h013c: oData <= 16'h0000;
            14'h013d: oData <= 16'h0000;
            14'h013e: oData <= 16'h0000;
            14'h013f: oData <= 16'h0000;
            14'h0140: oData <= 16'h02aa;
            14'h0141: oData <= 16'ha000;
            14'h0142: oData <= 16'h002a;
            14'h0143: oData <= 16'h02a8;
            14'h0144: oData <= 16'h0000;
            14'h0145: oData <= 16'hffe8;
            14'h0146: oData <= 16'hffff;
            14'h0147: oData <= 16'hfffb;
            14'h0148: oData <= 16'haaaf;
            14'h0149: oData <= 16'hfffe;
            14'h014a: oData <= 16'hfffe;
            14'h014b: oData <= 16'hfeff;
            14'h014c: oData <= 16'hffff;
            14'h014d: oData <= 16'hfeff;
            14'h014e: oData <= 16'habff;
            14'h014f: oData <= 16'h0000;
            14'h0150: oData <= 16'h0000;
            14'h0151: oData <= 16'h0000;
            14'h0152: oData <= 16'h0000;
            14'h0153: oData <= 16'h0000;
            14'h0154: oData <= 16'h0aaa;
            14'h0155: oData <= 16'ha000;
            14'h0156: oData <= 16'h00aa;
            14'h0157: oData <= 16'h02aa;
            14'h0158: oData <= 16'h0000;
            14'h0159: oData <= 16'hffea;
            14'h015a: oData <= 16'hffff;
            14'h015b: oData <= 16'hafff;
            14'h015c: oData <= 16'haaaa;
            14'h015d: oData <= 16'hffaa;
            14'h015e: oData <= 16'hfffe;
            14'h015f: oData <= 16'hfeff;
            14'h0160: oData <= 16'hffff;
            14'h0161: oData <= 16'hffff;
            14'h0162: oData <= 16'hafff;
            14'h0163: oData <= 16'h0000;
            14'h0164: oData <= 16'h0000;
            14'h0165: oData <= 16'h0000;
            14'h0166: oData <= 16'h0000;
            14'h0167: oData <= 16'h0000;
            14'h0168: oData <= 16'h0aa8;
            14'h0169: oData <= 16'h8000;
            14'h016a: oData <= 16'haaaa;
            14'h016b: oData <= 16'h02aa;
            14'h016c: oData <= 16'h8000;
            14'h016d: oData <= 16'hfffa;
            14'h016e: oData <= 16'hffff;
            14'h016f: oData <= 16'haaff;
            14'h0170: oData <= 16'heaaa;
            14'h0171: oData <= 16'hfaaa;
            14'h0172: oData <= 16'hffff;
            14'h0173: oData <= 16'hfeff;
            14'h0174: oData <= 16'hffff;
            14'h0175: oData <= 16'hffff;
            14'h0176: oData <= 16'hafff;
            14'h0177: oData <= 16'h0000;
            14'h0178: oData <= 16'h0000;
            14'h0179: oData <= 16'h0000;
            14'h017a: oData <= 16'h0000;
            14'h017b: oData <= 16'h0000;
            14'h017c: oData <= 16'h2aa8;
            14'h017d: oData <= 16'h0000;
            14'h017e: oData <= 16'haaaa;
            14'h017f: oData <= 16'h00aa;
            14'h0180: oData <= 16'ha000;
            14'h0181: oData <= 16'hfffe;
            14'h0182: oData <= 16'hffff;
            14'h0183: oData <= 16'haabf;
            14'h0184: oData <= 16'heaaa;
            14'h0185: oData <= 16'heabf;
            14'h0186: oData <= 16'hffff;
            14'h0187: oData <= 16'hfeff;
            14'h0188: oData <= 16'haaaa;
            14'h0189: oData <= 16'hfffa;
            14'h018a: oData <= 16'hafff;
            14'h018b: oData <= 16'h0002;
            14'h018c: oData <= 16'h0000;
            14'h018d: oData <= 16'h0000;
            14'h018e: oData <= 16'h0000;
            14'h018f: oData <= 16'h0000;
            14'h0190: oData <= 16'h2aa0;
            14'h0191: oData <= 16'h0000;
            14'h0192: oData <= 16'haaaa;
            14'h0193: oData <= 16'h00aa;
            14'h0194: oData <= 16'ha800;
            14'h0195: oData <= 16'hfaaa;
            14'h0196: oData <= 16'hafff;
            14'h0197: oData <= 16'hbeaf;
            14'h0198: oData <= 16'heaaa;
            14'h0199: oData <= 16'habff;
            14'h019a: oData <= 16'hfffe;
            14'h019b: oData <= 16'hafff;
            14'h019c: oData <= 16'hffaa;
            14'h019d: oData <= 16'hffab;
            14'h019e: oData <= 16'hbfff;
            14'h019f: oData <= 16'h002a;
            14'h01a0: oData <= 16'h0000;
            14'h01a1: oData <= 16'h0000;
            14'h01a2: oData <= 16'h0000;
            14'h01a3: oData <= 16'h0000;
            14'h01a4: oData <= 16'h2aa0;
            14'h01a5: oData <= 16'h0000;
            14'h01a6: oData <= 16'haaa8;
            14'h01a7: oData <= 16'h002a;
            14'h01a8: oData <= 16'haa00;
            14'h01a9: oData <= 16'hffff;
            14'h01aa: oData <= 16'hfaff;
            14'h01ab: oData <= 16'haaab;
            14'h01ac: oData <= 16'haaaa;
            14'h01ad: oData <= 16'haffe;
            14'h01ae: oData <= 16'hfffe;
            14'h01af: oData <= 16'habff;
            14'h01b0: oData <= 16'haaaa;
            14'h01b1: oData <= 16'hefaa;
            14'h01b2: oData <= 16'hffff;
            14'h01b3: oData <= 16'h00aa;
            14'h01b4: oData <= 16'h0000;
            14'h01b5: oData <= 16'h0000;
            14'h01b6: oData <= 16'h0000;
            14'h01b7: oData <= 16'h0000;
            14'h01b8: oData <= 16'haaa0;
            14'h01b9: oData <= 16'h0000;
            14'h01ba: oData <= 16'h0000;
            14'h01bb: oData <= 16'h0000;
            14'h01bc: oData <= 16'hba80;
            14'h01bd: oData <= 16'haaaa;
            14'h01be: oData <= 16'hebff;
            14'h01bf: oData <= 16'haaab;
            14'h01c0: oData <= 16'haaaa;
            14'h01c1: oData <= 16'hbfea;
            14'h01c2: oData <= 16'hfffa;
            14'h01c3: oData <= 16'haaeb;
            14'h01c4: oData <= 16'haaaa;
            14'h01c5: oData <= 16'habaa;
            14'h01c6: oData <= 16'heaab;
            14'h01c7: oData <= 16'h02af;
            14'h01c8: oData <= 16'h0000;
            14'h01c9: oData <= 16'h0000;
            14'h01ca: oData <= 16'h0000;
            14'h01cb: oData <= 16'h0000;
            14'h01cc: oData <= 16'haa80;
            14'h01cd: oData <= 16'h0000;
            14'h01ce: oData <= 16'h0000;
            14'h01cf: oData <= 16'h0000;
            14'h01d0: oData <= 16'heea0;
            14'h01d1: oData <= 16'hffff;
            14'h01d2: oData <= 16'hbfff;
            14'h01d3: oData <= 16'hfebe;
            14'h01d4: oData <= 16'hffff;
            14'h01d5: oData <= 16'haaaa;
            14'h01d6: oData <= 16'hfffe;
            14'h01d7: oData <= 16'haaaa;
            14'h01d8: oData <= 16'hfeaa;
            14'h01d9: oData <= 16'hffff;
            14'h01da: oData <= 16'hbffe;
            14'h01db: oData <= 16'h02bf;
            14'h01dc: oData <= 16'h0000;
            14'h01dd: oData <= 16'h0000;
            14'h01de: oData <= 16'h0000;
            14'h01df: oData <= 16'h0000;
            14'h01e0: oData <= 16'haa80;
            14'h01e1: oData <= 16'ha000;
            14'h01e2: oData <= 16'h0002;
            14'h01e3: oData <= 16'h0000;
            14'h01e4: oData <= 16'hfba8;
            14'h01e5: oData <= 16'haabf;
            14'h01e6: oData <= 16'hbfea;
            14'h01e7: oData <= 16'hffff;
            14'h01e8: oData <= 16'hfeaf;
            14'h01e9: oData <= 16'haaaf;
            14'h01ea: oData <= 16'hfffe;
            14'h01eb: oData <= 16'haaaf;
            14'h01ec: oData <= 16'hffff;
            14'h01ed: oData <= 16'hffff;
            14'h01ee: oData <= 16'hfaff;
            14'h01ef: oData <= 16'h0abe;
            14'h01f0: oData <= 16'h0000;
            14'h01f1: oData <= 16'h0000;
            14'h01f2: oData <= 16'h0000;
            14'h01f3: oData <= 16'h0000;
            14'h01f4: oData <= 16'haa80;
            14'h01f5: oData <= 16'ha802;
            14'h01f6: oData <= 16'h000a;
            14'h01f7: oData <= 16'h0000;
            14'h01f8: oData <= 16'hfeea;
            14'h01f9: oData <= 16'haaab;
            14'h01fa: oData <= 16'hfaaa;
            14'h01fb: oData <= 16'hffff;
            14'h01fc: oData <= 16'hffab;
            14'h01fd: oData <= 16'hebff;
            14'h01fe: oData <= 16'hffff;
            14'h01ff: oData <= 16'hfaff;
            14'h0200: oData <= 16'hffff;
            14'h0201: oData <= 16'hffff;
            14'h0202: oData <= 16'hefff;
            14'h0203: oData <= 16'h0aeb;
            14'h0204: oData <= 16'h0000;
            14'h0205: oData <= 16'h0000;
            14'h0206: oData <= 16'h0000;
            14'h0207: oData <= 16'h0000;
            14'h0208: oData <= 16'haa00;
            14'h0209: oData <= 16'haa82;
            14'h020a: oData <= 16'h000a;
            14'h020b: oData <= 16'h0000;
            14'h020c: oData <= 16'hffba;
            14'h020d: oData <= 16'hffaa;
            14'h020e: oData <= 16'haaaf;
            14'h020f: oData <= 16'hbfff;
            14'h0210: oData <= 16'hffea;
            14'h0211: oData <= 16'hffff;
            14'h0212: oData <= 16'hffff;
            14'h0213: oData <= 16'hfaff;
            14'h0214: oData <= 16'hffff;
            14'h0215: oData <= 16'hafff;
            14'h0216: oData <= 16'hbfaa;
            14'h0217: oData <= 16'h0aef;
            14'h0218: oData <= 16'h0000;
            14'h0219: oData <= 16'h0000;
            14'h021a: oData <= 16'h0000;
            14'h021b: oData <= 16'h0000;
            14'h021c: oData <= 16'haa00;
            14'h021d: oData <= 16'haaaa;
            14'h021e: oData <= 16'h000a;
            14'h021f: oData <= 16'h8000;
            14'h0220: oData <= 16'hffba;
            14'h0221: oData <= 16'hfffa;
            14'h0222: oData <= 16'haafe;
            14'h0223: oData <= 16'haaaa;
            14'h0224: oData <= 16'hfffa;
            14'h0225: oData <= 16'hffff;
            14'h0226: oData <= 16'hffff;
            14'h0227: oData <= 16'hfaff;
            14'h0228: oData <= 16'hffff;
            14'h0229: oData <= 16'habff;
            14'h022a: oData <= 16'hbaaa;
            14'h022b: oData <= 16'h0abf;
            14'h022c: oData <= 16'h0000;
            14'h022d: oData <= 16'h0000;
            14'h022e: oData <= 16'h0000;
            14'h022f: oData <= 16'h0000;
            14'h0230: oData <= 16'haa00;
            14'h0231: oData <= 16'haaaa;
            14'h0232: oData <= 16'h0002;
            14'h0233: oData <= 16'h8000;
            14'h0234: oData <= 16'hbfbe;
            14'h0235: oData <= 16'hbffa;
            14'h0236: oData <= 16'hbffe;
            14'h0237: oData <= 16'haaaa;
            14'h0238: oData <= 16'hffff;
            14'h0239: oData <= 16'hffff;
            14'h023a: oData <= 16'hffff;
            14'h023b: oData <= 16'hfaff;
            14'h023c: oData <= 16'hafff;
            14'h023d: oData <= 16'heabf;
            14'h023e: oData <= 16'hbabf;
            14'h023f: oData <= 16'h0abf;
            14'h0240: oData <= 16'h0000;
            14'h0241: oData <= 16'h0000;
            14'h0242: oData <= 16'h0000;
            14'h0243: oData <= 16'h0000;
            14'h0244: oData <= 16'ha800;
            14'h0245: oData <= 16'haaaa;
            14'h0246: oData <= 16'h0000;
            14'h0247: oData <= 16'ha000;
            14'h0248: oData <= 16'hbfbe;
            14'h0249: oData <= 16'hbffe;
            14'h024a: oData <= 16'hfffe;
            14'h024b: oData <= 16'hffff;
            14'h024c: oData <= 16'hffff;
            14'h024d: oData <= 16'hffff;
            14'h024e: oData <= 16'hffff;
            14'h024f: oData <= 16'hfaff;
            14'h0250: oData <= 16'hafff;
            14'h0251: oData <= 16'hfaaa;
            14'h0252: oData <= 16'hbbff;
            14'h0253: oData <= 16'h0abf;
            14'h0254: oData <= 16'h0000;
            14'h0255: oData <= 16'h0000;
            14'h0256: oData <= 16'h0000;
            14'h0257: oData <= 16'h0000;
            14'h0258: oData <= 16'ha800;
            14'h0259: oData <= 16'h0aaa;
            14'h025a: oData <= 16'h0000;
            14'h025b: oData <= 16'ha000;
            14'h025c: oData <= 16'hafbf;
            14'h025d: oData <= 16'hbffe;
            14'h025e: oData <= 16'hffea;
            14'h025f: oData <= 16'hffff;
            14'h0260: oData <= 16'hffff;
            14'h0261: oData <= 16'hffff;
            14'h0262: oData <= 16'hffff;
            14'h0263: oData <= 16'haaff;
            14'h0264: oData <= 16'hbfff;
            14'h0265: oData <= 16'hfeaa;
            14'h0266: oData <= 16'hfffe;
            14'h0267: oData <= 16'h0abe;
            14'h0268: oData <= 16'h0000;
            14'h0269: oData <= 16'h0000;
            14'h026a: oData <= 16'h0000;
            14'h026b: oData <= 16'h0000;
            14'h026c: oData <= 16'ha800;
            14'h026d: oData <= 16'h00aa;
            14'h026e: oData <= 16'h0000;
            14'h026f: oData <= 16'ha000;
            14'h0270: oData <= 16'hafbf;
            14'h0271: oData <= 16'hafff;
            14'h0272: oData <= 16'hfeaa;
            14'h0273: oData <= 16'hffff;
            14'h0274: oData <= 16'hffff;
            14'h0275: oData <= 16'haafb;
            14'h0276: oData <= 16'hffff;
            14'h0277: oData <= 16'habff;
            14'h0278: oData <= 16'hfffe;
            14'h0279: oData <= 16'hbfff;
            14'h027a: oData <= 16'hfffe;
            14'h027b: oData <= 16'h0abe;
            14'h027c: oData <= 16'h0000;
            14'h027d: oData <= 16'h0000;
            14'h027e: oData <= 16'h0000;
            14'h027f: oData <= 16'h0000;
            14'h0280: oData <= 16'ha000;
            14'h0281: oData <= 16'h000a;
            14'h0282: oData <= 16'h0000;
            14'h0283: oData <= 16'ha000;
            14'h0284: oData <= 16'hafbf;
            14'h0285: oData <= 16'haaff;
            14'h0286: oData <= 16'heaaf;
            14'h0287: oData <= 16'hffff;
            14'h0288: oData <= 16'hffff;
            14'h0289: oData <= 16'haabb;
            14'h028a: oData <= 16'hfffe;
            14'h028b: oData <= 16'hbfff;
            14'h028c: oData <= 16'hffea;
            14'h028d: oData <= 16'hbfff;
            14'h028e: oData <= 16'hfffe;
            14'h028f: oData <= 16'h0abe;
            14'h0290: oData <= 16'h0000;
            14'h0291: oData <= 16'h0000;
            14'h0292: oData <= 16'h0000;
            14'h0293: oData <= 16'h0000;
            14'h0294: oData <= 16'h0000;
            14'h0295: oData <= 16'h0000;
            14'h0296: oData <= 16'h0000;
            14'h0297: oData <= 16'ha000;
            14'h0298: oData <= 16'hafbe;
            14'h0299: oData <= 16'haaaf;
            14'h029a: oData <= 16'haaff;
            14'h029b: oData <= 16'hfffe;
            14'h029c: oData <= 16'haaab;
            14'h029d: oData <= 16'hfeae;
            14'h029e: oData <= 16'hffff;
            14'h029f: oData <= 16'hffff;
            14'h02a0: oData <= 16'hffaa;
            14'h02a1: oData <= 16'hbfff;
            14'h02a2: oData <= 16'hbffe;
            14'h02a3: oData <= 16'h0aef;
            14'h02a4: oData <= 16'h0000;
            14'h02a5: oData <= 16'h0000;
            14'h02a6: oData <= 16'h0000;
            14'h02a7: oData <= 16'h0000;
            14'h02a8: oData <= 16'h0000;
            14'h02a9: oData <= 16'h0000;
            14'h02aa: oData <= 16'h0000;
            14'h02ab: oData <= 16'h8000;
            14'h02ac: oData <= 16'hafbe;
            14'h02ad: oData <= 16'haeae;
            14'h02ae: oData <= 16'haffe;
            14'h02af: oData <= 16'hffaa;
            14'h02b0: oData <= 16'hfffb;
            14'h02b1: oData <= 16'hffaf;
            14'h02b2: oData <= 16'hffff;
            14'h02b3: oData <= 16'hffff;
            14'h02b4: oData <= 16'hfeaa;
            14'h02b5: oData <= 16'hbfff;
            14'h02b6: oData <= 16'hebea;
            14'h02b7: oData <= 16'h0aaf;
            14'h02b8: oData <= 16'h0000;
            14'h02b9: oData <= 16'h0000;
            14'h02ba: oData <= 16'h0000;
            14'h02bb: oData <= 16'h0000;
            14'h02bc: oData <= 16'h0000;
            14'h02bd: oData <= 16'h0000;
            14'h02be: oData <= 16'h0000;
            14'h02bf: oData <= 16'h8000;
            14'h02c0: oData <= 16'hbfbe;
            14'h02c1: oData <= 16'hbffe;
            14'h02c2: oData <= 16'hfffe;
            14'h02c3: oData <= 16'hfaaa;
            14'h02c4: oData <= 16'hffff;
            14'h02c5: oData <= 16'hbfaf;
            14'h02c6: oData <= 16'hfaaa;
            14'h02c7: oData <= 16'hbfff;
            14'h02c8: oData <= 16'hebaa;
            14'h02c9: oData <= 16'hbfff;
            14'h02ca: oData <= 16'hffea;
            14'h02cb: oData <= 16'h02bb;
            14'h02cc: oData <= 16'h0000;
            14'h02cd: oData <= 16'h0000;
            14'h02ce: oData <= 16'h0000;
            14'h02cf: oData <= 16'h0000;
            14'h02d0: oData <= 16'h0000;
            14'h02d1: oData <= 16'h0000;
            14'h02d2: oData <= 16'h0000;
            14'h02d3: oData <= 16'h8000;
            14'h02d4: oData <= 16'hbefe;
            14'h02d5: oData <= 16'hbffa;
            14'h02d6: oData <= 16'hfffa;
            14'h02d7: oData <= 16'haaaf;
            14'h02d8: oData <= 16'hfffe;
            14'h02d9: oData <= 16'hbeaf;
            14'h02da: oData <= 16'hfaaa;
            14'h02db: oData <= 16'hbfff;
            14'h02dc: oData <= 16'hbfae;
            14'h02dd: oData <= 16'haffe;
            14'h02de: oData <= 16'hafea;
            14'h02df: oData <= 16'h02be;
            14'h02e0: oData <= 16'h0000;
            14'h02e1: oData <= 16'h0000;
            14'h02e2: oData <= 16'h0000;
            14'h02e3: oData <= 16'h0000;
            14'h02e4: oData <= 16'h0000;
            14'h02e5: oData <= 16'h0000;
            14'h02e6: oData <= 16'h0000;
            14'h02e7: oData <= 16'h8000;
            14'h02e8: oData <= 16'hfefa;
            14'h02e9: oData <= 16'hbffa;
            14'h02ea: oData <= 16'hffea;
            14'h02eb: oData <= 16'habaf;
            14'h02ec: oData <= 16'hfeaa;
            14'h02ed: oData <= 16'hbabf;
            14'h02ee: oData <= 16'hffff;
            14'h02ef: oData <= 16'hafff;
            14'h02f0: oData <= 16'hfffe;
            14'h02f1: oData <= 16'habfb;
            14'h02f2: oData <= 16'hfbeb;
            14'h02f3: oData <= 16'h02af;
            14'h02f4: oData <= 16'h0000;
            14'h02f5: oData <= 16'h0000;
            14'h02f6: oData <= 16'h0000;
            14'h02f7: oData <= 16'h0000;
            14'h02f8: oData <= 16'h0000;
            14'h02f9: oData <= 16'h0000;
            14'h02fa: oData <= 16'h0000;
            14'h02fb: oData <= 16'h0000;
            14'h02fc: oData <= 16'hfbea;
            14'h02fd: oData <= 16'hbfff;
            14'h02fe: oData <= 16'hfeaa;
            14'h02ff: oData <= 16'hffaf;
            14'h0300: oData <= 16'haaaa;
            14'h0301: oData <= 16'hfeff;
            14'h0302: oData <= 16'hffff;
            14'h0303: oData <= 16'haaeb;
            14'h0304: oData <= 16'hffff;
            14'h0305: oData <= 16'haaff;
            14'h0306: oData <= 16'hffea;
            14'h0307: oData <= 16'h00ab;
            14'h0308: oData <= 16'h0000;
            14'h0309: oData <= 16'h0000;
            14'h030a: oData <= 16'h0000;
            14'h030b: oData <= 16'h0000;
            14'h030c: oData <= 16'h0000;
            14'h030d: oData <= 16'h0000;
            14'h030e: oData <= 16'h0000;
            14'h030f: oData <= 16'h0000;
            14'h0310: oData <= 16'hafe8;
            14'h0311: oData <= 16'hffff;
            14'h0312: oData <= 16'heaaa;
            14'h0313: oData <= 16'hffaf;
            14'h0314: oData <= 16'haaff;
            14'h0315: oData <= 16'hffea;
            14'h0316: oData <= 16'hffff;
            14'h0317: oData <= 16'heaab;
            14'h0318: oData <= 16'hffff;
            14'h0319: oData <= 16'hbaaf;
            14'h031a: oData <= 16'hffaa;
            14'h031b: oData <= 16'h002b;
            14'h031c: oData <= 16'h0000;
            14'h031d: oData <= 16'h0000;
            14'h031e: oData <= 16'h0000;
            14'h031f: oData <= 16'h0000;
            14'h0320: oData <= 16'h0000;
            14'h0321: oData <= 16'h0000;
            14'h0322: oData <= 16'h0000;
            14'h0323: oData <= 16'h0000;
            14'h0324: oData <= 16'hffa8;
            14'h0325: oData <= 16'hfffa;
            14'h0326: oData <= 16'haaab;
            14'h0327: oData <= 16'hfeae;
            14'h0328: oData <= 16'hbfff;
            14'h0329: oData <= 16'heaaa;
            14'h032a: oData <= 16'hffff;
            14'h032b: oData <= 16'hfeaf;
            14'h032c: oData <= 16'hffff;
            14'h032d: oData <= 16'hbaaa;
            14'h032e: oData <= 16'hffae;
            14'h032f: oData <= 16'h002a;
            14'h0330: oData <= 16'h0000;
            14'h0331: oData <= 16'h0000;
            14'h0332: oData <= 16'h0000;
            14'h0333: oData <= 16'h0000;
            14'h0334: oData <= 16'h0000;
            14'h0335: oData <= 16'h0000;
            14'h0336: oData <= 16'h0000;
            14'h0337: oData <= 16'h0000;
            14'h0338: oData <= 16'heaa0;
            14'h0339: oData <= 16'hffff;
            14'h033a: oData <= 16'habaf;
            14'h033b: oData <= 16'hfaaa;
            14'h033c: oData <= 16'hffff;
            14'h033d: oData <= 16'haaaa;
            14'h033e: oData <= 16'hfeaa;
            14'h033f: oData <= 16'hffff;
            14'h0340: oData <= 16'habff;
            14'h0341: oData <= 16'hbaea;
            14'h0342: oData <= 16'hffaa;
            14'h0343: oData <= 16'h000a;
            14'h0344: oData <= 16'h0000;
            14'h0345: oData <= 16'h0000;
            14'h0346: oData <= 16'h0000;
            14'h0347: oData <= 16'h0000;
            14'h0348: oData <= 16'h0000;
            14'h0349: oData <= 16'h0000;
            14'h034a: oData <= 16'h0000;
            14'h034b: oData <= 16'h0000;
            14'h034c: oData <= 16'hba80;
            14'h034d: oData <= 16'hffff;
            14'h034e: oData <= 16'hfeaf;
            14'h034f: oData <= 16'heaaa;
            14'h0350: oData <= 16'hffff;
            14'h0351: oData <= 16'haffa;
            14'h0352: oData <= 16'haaaa;
            14'h0353: oData <= 16'haaaa;
            14'h0354: oData <= 16'haaaa;
            14'h0355: oData <= 16'hfafe;
            14'h0356: oData <= 16'hffaa;
            14'h0357: oData <= 16'h000a;
            14'h0358: oData <= 16'h0000;
            14'h0359: oData <= 16'h0000;
            14'h035a: oData <= 16'h0000;
            14'h035b: oData <= 16'h0000;
            14'h035c: oData <= 16'h0000;
            14'h035d: oData <= 16'h0000;
            14'h035e: oData <= 16'h0000;
            14'h035f: oData <= 16'h0000;
            14'h0360: oData <= 16'hea00;
            14'h0361: oData <= 16'hffff;
            14'h0362: oData <= 16'hfabf;
            14'h0363: oData <= 16'haaaf;
            14'h0364: oData <= 16'hfffa;
            14'h0365: oData <= 16'hfffa;
            14'h0366: oData <= 16'haaff;
            14'h0367: oData <= 16'haaaa;
            14'h0368: oData <= 16'haaaa;
            14'h0369: oData <= 16'hfaff;
            14'h036a: oData <= 16'hffaa;
            14'h036b: oData <= 16'h000a;
            14'h036c: oData <= 16'h0000;
            14'h036d: oData <= 16'h0000;
            14'h036e: oData <= 16'h0000;
            14'h036f: oData <= 16'h0000;
            14'h0370: oData <= 16'h0000;
            14'h0371: oData <= 16'h0000;
            14'h0372: oData <= 16'h0000;
            14'h0373: oData <= 16'h0000;
            14'h0374: oData <= 16'ha800;
            14'h0375: oData <= 16'hffff;
            14'h0376: oData <= 16'hfaff;
            14'h0377: oData <= 16'haaaf;
            14'h0378: oData <= 16'hbeaa;
            14'h0379: oData <= 16'hfffa;
            14'h037a: oData <= 16'hfaff;
            14'h037b: oData <= 16'hebff;
            14'h037c: oData <= 16'hafff;
            14'h037d: oData <= 16'hfafe;
            14'h037e: oData <= 16'hffaa;
            14'h037f: oData <= 16'h000a;
            14'h0380: oData <= 16'h0000;
            14'h0381: oData <= 16'h0000;
            14'h0382: oData <= 16'h0000;
            14'h0383: oData <= 16'h0000;
            14'h0384: oData <= 16'h0000;
            14'h0385: oData <= 16'h0000;
            14'h0386: oData <= 16'h0000;
            14'h0387: oData <= 16'h0000;
            14'h0388: oData <= 16'ha000;
            14'h0389: oData <= 16'hfffe;
            14'h038a: oData <= 16'heaff;
            14'h038b: oData <= 16'hafaf;
            14'h038c: oData <= 16'haaaa;
            14'h038d: oData <= 16'hfffe;
            14'h038e: oData <= 16'hfaff;
            14'h038f: oData <= 16'hebff;
            14'h0390: oData <= 16'hbfff;
            14'h0391: oData <= 16'hbafe;
            14'h0392: oData <= 16'hffaa;
            14'h0393: oData <= 16'h000a;
            14'h0394: oData <= 16'h0000;
            14'h0395: oData <= 16'h0000;
            14'h0396: oData <= 16'h0000;
            14'h0397: oData <= 16'h0000;
            14'h0398: oData <= 16'h0000;
            14'h0399: oData <= 16'h0000;
            14'h039a: oData <= 16'h0000;
            14'h039b: oData <= 16'h0000;
            14'h039c: oData <= 16'h8000;
            14'h039d: oData <= 16'hfffa;
            14'h039e: oData <= 16'habff;
            14'h039f: oData <= 16'hffaf;
            14'h03a0: oData <= 16'haaaa;
            14'h03a1: oData <= 16'hffea;
            14'h03a2: oData <= 16'hfaff;
            14'h03a3: oData <= 16'hebff;
            14'h03a4: oData <= 16'hbfff;
            14'h03a5: oData <= 16'haafe;
            14'h03a6: oData <= 16'hffaa;
            14'h03a7: oData <= 16'h000a;
            14'h03a8: oData <= 16'h0000;
            14'h03a9: oData <= 16'h0000;
            14'h03aa: oData <= 16'h0000;
            14'h03ab: oData <= 16'h0000;
            14'h03ac: oData <= 16'h0000;
            14'h03ad: oData <= 16'h0000;
            14'h03ae: oData <= 16'h0000;
            14'h03af: oData <= 16'h0000;
            14'h03b0: oData <= 16'h0000;
            14'h03b1: oData <= 16'hfffa;
            14'h03b2: oData <= 16'hafff;
            14'h03b3: oData <= 16'hffae;
            14'h03b4: oData <= 16'haaaf;
            14'h03b5: oData <= 16'heaaa;
            14'h03b6: oData <= 16'hfaff;
            14'h03b7: oData <= 16'hebff;
            14'h03b8: oData <= 16'haaff;
            14'h03b9: oData <= 16'haaaa;
            14'h03ba: oData <= 16'hffaa;
            14'h03bb: oData <= 16'h000a;
            14'h03bc: oData <= 16'h0000;
            14'h03bd: oData <= 16'h0000;
            14'h03be: oData <= 16'h0000;
            14'h03bf: oData <= 16'h0000;
            14'h03c0: oData <= 16'h0000;
            14'h03c1: oData <= 16'h0000;
            14'h03c2: oData <= 16'h0000;
            14'h03c3: oData <= 16'h0000;
            14'h03c4: oData <= 16'h0000;
            14'h03c5: oData <= 16'hfffa;
            14'h03c6: oData <= 16'hbfff;
            14'h03c7: oData <= 16'hffaa;
            14'h03c8: oData <= 16'hafff;
            14'h03c9: oData <= 16'haaaa;
            14'h03ca: oData <= 16'haaaa;
            14'h03cb: oData <= 16'haaaa;
            14'h03cc: oData <= 16'haaaa;
            14'h03cd: oData <= 16'haaaa;
            14'h03ce: oData <= 16'hffaa;
            14'h03cf: oData <= 16'h000a;
            14'h03d0: oData <= 16'h0000;
            14'h03d1: oData <= 16'h0000;
            14'h03d2: oData <= 16'h0000;
            14'h03d3: oData <= 16'h0000;
            14'h03d4: oData <= 16'h0000;
            14'h03d5: oData <= 16'h0000;
            14'h03d6: oData <= 16'h0000;
            14'h03d7: oData <= 16'h0000;
            14'h03d8: oData <= 16'h0000;
            14'h03d9: oData <= 16'hffea;
            14'h03da: oData <= 16'hffff;
            14'h03db: oData <= 16'hffea;
            14'h03dc: oData <= 16'hafff;
            14'h03dd: oData <= 16'haaab;
            14'h03de: oData <= 16'haaaa;
            14'h03df: oData <= 16'haaaa;
            14'h03e0: oData <= 16'haaaa;
            14'h03e1: oData <= 16'haaaa;
            14'h03e2: oData <= 16'hffaa;
            14'h03e3: oData <= 16'h000a;
            14'h03e4: oData <= 16'h0000;
            14'h03e5: oData <= 16'h0000;
            14'h03e6: oData <= 16'h0000;
            14'h03e7: oData <= 16'h0000;
            14'h03e8: oData <= 16'h0000;
            14'h03e9: oData <= 16'h0000;
            14'h03ea: oData <= 16'h0000;
            14'h03eb: oData <= 16'h0000;
            14'h03ec: oData <= 16'h0000;
            14'h03ed: oData <= 16'hffe8;
            14'h03ee: oData <= 16'hffff;
            14'h03ef: oData <= 16'hffab;
            14'h03f0: oData <= 16'hafff;
            14'h03f1: oData <= 16'haaff;
            14'h03f2: oData <= 16'haaaa;
            14'h03f3: oData <= 16'haaaa;
            14'h03f4: oData <= 16'haaaa;
            14'h03f5: oData <= 16'haaaa;
            14'h03f6: oData <= 16'hffaa;
            14'h03f7: oData <= 16'h000a;
            14'h03f8: oData <= 16'h0000;
            14'h03f9: oData <= 16'h0000;
            14'h03fa: oData <= 16'h0000;
            14'h03fb: oData <= 16'h0000;
            14'h03fc: oData <= 16'h0000;
            14'h03fd: oData <= 16'h0000;
            14'h03fe: oData <= 16'h0000;
            14'h03ff: oData <= 16'h0000;
            14'h0400: oData <= 16'h0000;
            14'h0401: oData <= 16'hffa8;
            14'h0402: oData <= 16'hffff;
            14'h0403: oData <= 16'hfeaf;
            14'h0404: oData <= 16'hafff;
            14'h0405: oData <= 16'hbfff;
            14'h0406: oData <= 16'haaaa;
            14'h0407: oData <= 16'haaaa;
            14'h0408: oData <= 16'haaaa;
            14'h0409: oData <= 16'haaaa;
            14'h040a: oData <= 16'hffea;
            14'h040b: oData <= 16'h000a;
            14'h040c: oData <= 16'h0000;
            14'h040d: oData <= 16'h0000;
            14'h040e: oData <= 16'h0000;
            14'h040f: oData <= 16'h0000;
            14'h0410: oData <= 16'h0000;
            14'h0411: oData <= 16'h0000;
            14'h0412: oData <= 16'h0000;
            14'h0413: oData <= 16'h0000;
            14'h0414: oData <= 16'h0000;
            14'h0415: oData <= 16'hfea0;
            14'h0416: oData <= 16'hffff;
            14'h0417: oData <= 16'heabf;
            14'h0418: oData <= 16'habff;
            14'h0419: oData <= 16'hffff;
            14'h041a: oData <= 16'haaaf;
            14'h041b: oData <= 16'haaaa;
            14'h041c: oData <= 16'haaaa;
            14'h041d: oData <= 16'haaaa;
            14'h041e: oData <= 16'hffeb;
            14'h041f: oData <= 16'h000a;
            14'h0420: oData <= 16'h0000;
            14'h0421: oData <= 16'h0000;
            14'h0422: oData <= 16'h0000;
            14'h0423: oData <= 16'h0000;
            14'h0424: oData <= 16'h0000;
            14'h0425: oData <= 16'h0000;
            14'h0426: oData <= 16'h0000;
            14'h0427: oData <= 16'h0000;
            14'h0428: oData <= 16'h0000;
            14'h0429: oData <= 16'hfa80;
            14'h042a: oData <= 16'hffff;
            14'h042b: oData <= 16'haaff;
            14'h042c: oData <= 16'hebff;
            14'h042d: oData <= 16'hffff;
            14'h042e: oData <= 16'hbfaf;
            14'h042f: oData <= 16'haaaa;
            14'h0430: oData <= 16'haaaa;
            14'h0431: oData <= 16'hafaa;
            14'h0432: oData <= 16'hffeb;
            14'h0433: oData <= 16'h000a;
            14'h0434: oData <= 16'h0000;
            14'h0435: oData <= 16'h0000;
            14'h0436: oData <= 16'h0000;
            14'h0437: oData <= 16'h0000;
            14'h0438: oData <= 16'h0000;
            14'h0439: oData <= 16'h0000;
            14'h043a: oData <= 16'h0000;
            14'h043b: oData <= 16'h0000;
            14'h043c: oData <= 16'h0000;
            14'h043d: oData <= 16'hea00;
            14'h043e: oData <= 16'hffff;
            14'h043f: oData <= 16'hafff;
            14'h0440: oData <= 16'hebfa;
            14'h0441: oData <= 16'hffff;
            14'h0442: oData <= 16'hffaf;
            14'h0443: oData <= 16'heaff;
            14'h0444: oData <= 16'hfaff;
            14'h0445: oData <= 16'hebeb;
            14'h0446: oData <= 16'hfffa;
            14'h0447: oData <= 16'h000a;
            14'h0448: oData <= 16'h0000;
            14'h0449: oData <= 16'h0000;
            14'h044a: oData <= 16'h0000;
            14'h044b: oData <= 16'h0000;
            14'h044c: oData <= 16'h0000;
            14'h044d: oData <= 16'h0000;
            14'h044e: oData <= 16'h0000;
            14'h044f: oData <= 16'h0000;
            14'h0450: oData <= 16'h0000;
            14'h0451: oData <= 16'haa00;
            14'h0452: oData <= 16'hffff;
            14'h0453: oData <= 16'hbfff;
            14'h0454: oData <= 16'heaaa;
            14'h0455: oData <= 16'hffff;
            14'h0456: oData <= 16'hffaf;
            14'h0457: oData <= 16'hfaff;
            14'h0458: oData <= 16'hfabf;
            14'h0459: oData <= 16'haaea;
            14'h045a: oData <= 16'hfffa;
            14'h045b: oData <= 16'h000a;
            14'h045c: oData <= 16'h0000;
            14'h045d: oData <= 16'h0000;
            14'h045e: oData <= 16'h0000;
            14'h045f: oData <= 16'h0000;
            14'h0460: oData <= 16'h0000;
            14'h0461: oData <= 16'h0000;
            14'h0462: oData <= 16'h0000;
            14'h0463: oData <= 16'h0000;
            14'h0464: oData <= 16'h0000;
            14'h0465: oData <= 16'ha000;
            14'h0466: oData <= 16'hffbe;
            14'h0467: oData <= 16'hfffa;
            14'h0468: oData <= 16'hfaab;
            14'h0469: oData <= 16'hffff;
            14'h046a: oData <= 16'hffaf;
            14'h046b: oData <= 16'hfaff;
            14'h046c: oData <= 16'hfebf;
            14'h046d: oData <= 16'hbbfa;
            14'h046e: oData <= 16'hfffe;
            14'h046f: oData <= 16'h000a;
            14'h0470: oData <= 16'h0000;
            14'h0471: oData <= 16'h0000;
            14'h0472: oData <= 16'h0000;
            14'h0473: oData <= 16'h0000;
            14'h0474: oData <= 16'h0000;
            14'h0475: oData <= 16'h0000;
            14'h0476: oData <= 16'h0000;
            14'h0477: oData <= 16'h0000;
            14'h0478: oData <= 16'h0000;
            14'h0479: oData <= 16'h8000;
            14'h047a: oData <= 16'hfafa;
            14'h047b: oData <= 16'hffbf;
            14'h047c: oData <= 16'haabf;
            14'h047d: oData <= 16'hfffe;
            14'h047e: oData <= 16'hffaf;
            14'h047f: oData <= 16'hfaff;
            14'h0480: oData <= 16'hbeaf;
            14'h0481: oData <= 16'haffa;
            14'h0482: oData <= 16'hfffe;
            14'h0483: oData <= 16'h000a;
            14'h0484: oData <= 16'h0000;
            14'h0485: oData <= 16'h0000;
            14'h0486: oData <= 16'h0000;
            14'h0487: oData <= 16'h0000;
            14'h0488: oData <= 16'h0000;
            14'h0489: oData <= 16'h0000;
            14'h048a: oData <= 16'h0000;
            14'h048b: oData <= 16'h0000;
            14'h048c: oData <= 16'h0000;
            14'h048d: oData <= 16'h0000;
            14'h048e: oData <= 16'hafea;
            14'h048f: oData <= 16'hfaff;
            14'h0490: oData <= 16'habff;
            14'h0491: oData <= 16'hffaa;
            14'h0492: oData <= 16'hffaf;
            14'h0493: oData <= 16'hfabf;
            14'h0494: oData <= 16'hffaf;
            14'h0495: oData <= 16'heaaa;
            14'h0496: oData <= 16'hffff;
            14'h0497: oData <= 16'h000a;
            14'h0498: oData <= 16'h0000;
            14'h0499: oData <= 16'h0000;
            14'h049a: oData <= 16'h0000;
            14'h049b: oData <= 16'h0000;
            14'h049c: oData <= 16'h0000;
            14'h049d: oData <= 16'h0000;
            14'h049e: oData <= 16'h0000;
            14'h049f: oData <= 16'h0000;
            14'h04a0: oData <= 16'h0000;
            14'h04a1: oData <= 16'h0000;
            14'h04a2: oData <= 16'hfea8;
            14'h04a3: oData <= 16'haffa;
            14'h04a4: oData <= 16'hffff;
            14'h04a5: oData <= 16'haaaa;
            14'h04a6: oData <= 16'hfeaa;
            14'h04a7: oData <= 16'hfebf;
            14'h04a8: oData <= 16'haaab;
            14'h04a9: oData <= 16'hfaaa;
            14'h04aa: oData <= 16'hffff;
            14'h04ab: oData <= 16'h000a;
            14'h04ac: oData <= 16'h0000;
            14'h04ad: oData <= 16'h0000;
            14'h04ae: oData <= 16'h0000;
            14'h04af: oData <= 16'h0000;
            14'h04b0: oData <= 16'h0000;
            14'h04b1: oData <= 16'h0000;
            14'h04b2: oData <= 16'h0000;
            14'h04b3: oData <= 16'h0000;
            14'h04b4: oData <= 16'h0000;
            14'h04b5: oData <= 16'h0000;
            14'h04b6: oData <= 16'hfaa0;
            14'h04b7: oData <= 16'hffaf;
            14'h04b8: oData <= 16'hfffa;
            14'h04b9: oData <= 16'haabf;
            14'h04ba: oData <= 16'haaaa;
            14'h04bb: oData <= 16'haaaa;
            14'h04bc: oData <= 16'haaaa;
            14'h04bd: oData <= 16'hfffa;
            14'h04be: oData <= 16'hffff;
            14'h04bf: oData <= 16'h000a;
            14'h04c0: oData <= 16'h0000;
            14'h04c1: oData <= 16'h0000;
            14'h04c2: oData <= 16'h0000;
            14'h04c3: oData <= 16'h0000;
            14'h04c4: oData <= 16'h0000;
            14'h04c5: oData <= 16'h0000;
            14'h04c6: oData <= 16'h0000;
            14'h04c7: oData <= 16'h0000;
            14'h04c8: oData <= 16'h0000;
            14'h04c9: oData <= 16'h0000;
            14'h04ca: oData <= 16'haa00;
            14'h04cb: oData <= 16'hfaff;
            14'h04cc: oData <= 16'hffaf;
            14'h04cd: oData <= 16'hffff;
            14'h04ce: oData <= 16'haaff;
            14'h04cf: oData <= 16'haaaa;
            14'h04d0: oData <= 16'hfffa;
            14'h04d1: oData <= 16'hffff;
            14'h04d2: oData <= 16'hffff;
            14'h04d3: oData <= 16'h000a;
            14'h04d4: oData <= 16'h0000;
            14'h04d5: oData <= 16'h0000;
            14'h04d6: oData <= 16'h0000;
            14'h04d7: oData <= 16'h0000;
            14'h04d8: oData <= 16'h0000;
            14'h04d9: oData <= 16'h0000;
            14'h04da: oData <= 16'h0000;
            14'h04db: oData <= 16'h0000;
            14'h04dc: oData <= 16'h0000;
            14'h04dd: oData <= 16'h0000;
            14'h04de: oData <= 16'ha800;
            14'h04df: oData <= 16'haffa;
            14'h04e0: oData <= 16'heaff;
            14'h04e1: oData <= 16'hffff;
            14'h04e2: oData <= 16'hffff;
            14'h04e3: oData <= 16'hffff;
            14'h04e4: oData <= 16'hffff;
            14'h04e5: oData <= 16'hbfff;
            14'h04e6: oData <= 16'hffff;
            14'h04e7: oData <= 16'h002a;
            14'h04e8: oData <= 16'h0000;
            14'h04e9: oData <= 16'h0000;
            14'h04ea: oData <= 16'h0000;
            14'h04eb: oData <= 16'h0000;
            14'h04ec: oData <= 16'h0000;
            14'h04ed: oData <= 16'h0000;
            14'h04ee: oData <= 16'h0000;
            14'h04ef: oData <= 16'h0000;
            14'h04f0: oData <= 16'h0000;
            14'h04f1: oData <= 16'h0000;
            14'h04f2: oData <= 16'h8000;
            14'h04f3: oData <= 16'hffaa;
            14'h04f4: oData <= 16'hbffa;
            14'h04f5: oData <= 16'hfffa;
            14'h04f6: oData <= 16'hffff;
            14'h04f7: oData <= 16'hffff;
            14'h04f8: oData <= 16'hffff;
            14'h04f9: oData <= 16'hefff;
            14'h04fa: oData <= 16'hffbf;
            14'h04fb: oData <= 16'h002b;
            14'h04fc: oData <= 16'h0000;
            14'h04fd: oData <= 16'h0000;
            14'h04fe: oData <= 16'h0000;
            14'h04ff: oData <= 16'h0000;
            14'h0500: oData <= 16'h0000;
            14'h0501: oData <= 16'h0000;
            14'h0502: oData <= 16'h0000;
            14'h0503: oData <= 16'h0000;
            14'h0504: oData <= 16'h0000;
            14'h0505: oData <= 16'h0000;
            14'h0506: oData <= 16'h0000;
            14'h0507: oData <= 16'hfaa8;
            14'h0508: oData <= 16'hfeaf;
            14'h0509: oData <= 16'hffaf;
            14'h050a: oData <= 16'haaff;
            14'h050b: oData <= 16'haaaa;
            14'h050c: oData <= 16'hffaa;
            14'h050d: oData <= 16'hfaff;
            14'h050e: oData <= 16'hffbf;
            14'h050f: oData <= 16'h002b;
            14'h0510: oData <= 16'h0000;
            14'h0511: oData <= 16'h0000;
            14'h0512: oData <= 16'h0000;
            14'h0513: oData <= 16'h0000;
            14'h0514: oData <= 16'h0000;
            14'h0515: oData <= 16'h0000;
            14'h0516: oData <= 16'h0000;
            14'h0517: oData <= 16'h0000;
            14'h0518: oData <= 16'h0000;
            14'h0519: oData <= 16'h0000;
            14'h051a: oData <= 16'h0000;
            14'h051b: oData <= 16'haa80;
            14'h051c: oData <= 16'habff;
            14'h051d: oData <= 16'haaff;
            14'h051e: oData <= 16'hfffe;
            14'h051f: oData <= 16'hffff;
            14'h0520: oData <= 16'hffff;
            14'h0521: oData <= 16'hffbf;
            14'h0522: oData <= 16'hffbf;
            14'h0523: oData <= 16'h002b;
            14'h0524: oData <= 16'h0000;
            14'h0525: oData <= 16'h0000;
            14'h0526: oData <= 16'h0000;
            14'h0527: oData <= 16'h0000;
            14'h0528: oData <= 16'h0000;
            14'h0529: oData <= 16'h0000;
            14'h052a: oData <= 16'h0000;
            14'h052b: oData <= 16'h0000;
            14'h052c: oData <= 16'h0000;
            14'h052d: oData <= 16'h0000;
            14'h052e: oData <= 16'h0000;
            14'h052f: oData <= 16'ha800;
            14'h0530: oData <= 16'hffea;
            14'h0531: oData <= 16'hffea;
            14'h0532: oData <= 16'haaab;
            14'h0533: oData <= 16'hffaa;
            14'h0534: oData <= 16'hbfff;
            14'h0535: oData <= 16'hffea;
            14'h0536: oData <= 16'hffef;
            14'h0537: oData <= 16'h002b;
            14'h0538: oData <= 16'h0000;
            14'h0539: oData <= 16'h0000;
            14'h053a: oData <= 16'h0000;
            14'h053b: oData <= 16'h0000;
            14'h053c: oData <= 16'h0000;
            14'h053d: oData <= 16'h0000;
            14'h053e: oData <= 16'h0000;
            14'h053f: oData <= 16'h0000;
            14'h0540: oData <= 16'ha000;
            14'h0541: oData <= 16'h0002;
            14'h0542: oData <= 16'h0000;
            14'h0543: oData <= 16'h8000;
            14'h0544: oData <= 16'hfeaa;
            14'h0545: oData <= 16'haabf;
            14'h0546: oData <= 16'hffff;
            14'h0547: oData <= 16'haaff;
            14'h0548: oData <= 16'heaaa;
            14'h0549: oData <= 16'hffff;
            14'h054a: oData <= 16'hfffa;
            14'h054b: oData <= 16'h002b;
            14'h054c: oData <= 16'h0000;
            14'h054d: oData <= 16'h0000;
            14'h054e: oData <= 16'h0000;
            14'h054f: oData <= 16'h0000;
            14'h0550: oData <= 16'h0000;
            14'h0551: oData <= 16'h0000;
            14'h0552: oData <= 16'h0000;
            14'h0553: oData <= 16'h0000;
            14'h0554: oData <= 16'ha800;
            14'h0555: oData <= 16'h000a;
            14'h0556: oData <= 16'h0000;
            14'h0557: oData <= 16'h0000;
            14'h0558: oData <= 16'heaa0;
            14'h0559: oData <= 16'hffff;
            14'h055a: oData <= 16'hfaaa;
            14'h055b: oData <= 16'hffff;
            14'h055c: oData <= 16'hffff;
            14'h055d: oData <= 16'hbfff;
            14'h055e: oData <= 16'hffff;
            14'h055f: oData <= 16'h002b;
            14'h0560: oData <= 16'h0000;
            14'h0561: oData <= 16'h0000;
            14'h0562: oData <= 16'h0000;
            14'h0563: oData <= 16'h0000;
            14'h0564: oData <= 16'h0000;
            14'h0565: oData <= 16'h0000;
            14'h0566: oData <= 16'h0000;
            14'h0567: oData <= 16'h0000;
            14'h0568: oData <= 16'ha800;
            14'h0569: oData <= 16'h000a;
            14'h056a: oData <= 16'h0000;
            14'h056b: oData <= 16'h0000;
            14'h056c: oData <= 16'haa00;
            14'h056d: oData <= 16'hfffe;
            14'h056e: oData <= 16'hafff;
            14'h056f: oData <= 16'haaaa;
            14'h0570: oData <= 16'hffff;
            14'h0571: oData <= 16'heabf;
            14'h0572: oData <= 16'hffff;
            14'h0573: oData <= 16'h002a;
            14'h0574: oData <= 16'h0000;
            14'h0575: oData <= 16'h0000;
            14'h0576: oData <= 16'h0000;
            14'h0577: oData <= 16'h0000;
            14'h0578: oData <= 16'h0000;
            14'h0579: oData <= 16'h0000;
            14'h057a: oData <= 16'h0000;
            14'h057b: oData <= 16'h0000;
            14'h057c: oData <= 16'ha800;
            14'h057d: oData <= 16'h002a;
            14'h057e: oData <= 16'h0000;
            14'h057f: oData <= 16'h0000;
            14'h0580: oData <= 16'ha000;
            14'h0581: oData <= 16'hffaa;
            14'h0582: oData <= 16'hffff;
            14'h0583: oData <= 16'hffff;
            14'h0584: oData <= 16'haaaa;
            14'h0585: oData <= 16'hffea;
            14'h0586: oData <= 16'hffff;
            14'h0587: oData <= 16'h000a;
            14'h0588: oData <= 16'h0a80;
            14'h0589: oData <= 16'h0000;
            14'h058a: oData <= 16'h0000;
            14'h058b: oData <= 16'h0000;
            14'h058c: oData <= 16'h0000;
            14'h058d: oData <= 16'h0000;
            14'h058e: oData <= 16'h0000;
            14'h058f: oData <= 16'h0000;
            14'h0590: oData <= 16'ha000;
            14'h0591: oData <= 16'h00aa;
            14'h0592: oData <= 16'h0000;
            14'h0593: oData <= 16'h0000;
            14'h0594: oData <= 16'h0000;
            14'h0595: oData <= 16'hfeaa;
            14'h0596: oData <= 16'hffff;
            14'h0597: oData <= 16'hffff;
            14'h0598: oData <= 16'hffff;
            14'h0599: oData <= 16'hffff;
            14'h059a: oData <= 16'hbfff;
            14'h059b: oData <= 16'h000a;
            14'h059c: oData <= 16'h2aa0;
            14'h059d: oData <= 16'h0000;
            14'h059e: oData <= 16'h0000;
            14'h059f: oData <= 16'h0000;
            14'h05a0: oData <= 16'h0000;
            14'h05a1: oData <= 16'h0000;
            14'h05a2: oData <= 16'h0000;
            14'h05a3: oData <= 16'h0000;
            14'h05a4: oData <= 16'h8000;
            14'h05a5: oData <= 16'h02aa;
            14'h05a6: oData <= 16'h0000;
            14'h05a7: oData <= 16'h0000;
            14'h05a8: oData <= 16'h0000;
            14'h05a9: oData <= 16'heaaa;
            14'h05aa: oData <= 16'hffff;
            14'h05ab: oData <= 16'hffff;
            14'h05ac: oData <= 16'hffff;
            14'h05ad: oData <= 16'hffff;
            14'h05ae: oData <= 16'hbfff;
            14'h05af: oData <= 16'h0002;
            14'h05b0: oData <= 16'h2aa8;
            14'h05b1: oData <= 16'h0000;
            14'h05b2: oData <= 16'h0000;
            14'h05b3: oData <= 16'h0000;
            14'h05b4: oData <= 16'h0000;
            14'h05b5: oData <= 16'h0000;
            14'h05b6: oData <= 16'h0000;
            14'h05b7: oData <= 16'h0000;
            14'h05b8: oData <= 16'h0000;
            14'h05b9: oData <= 16'h0aaa;
            14'h05ba: oData <= 16'h0000;
            14'h05bb: oData <= 16'h0000;
            14'h05bc: oData <= 16'h0000;
            14'h05bd: oData <= 16'haaaa;
            14'h05be: oData <= 16'hffaa;
            14'h05bf: oData <= 16'hffff;
            14'h05c0: oData <= 16'hffff;
            14'h05c1: oData <= 16'hffff;
            14'h05c2: oData <= 16'hafff;
            14'h05c3: oData <= 16'h0002;
            14'h05c4: oData <= 16'h0aa8;
            14'h05c5: oData <= 16'h0000;
            14'h05c6: oData <= 16'h0000;
            14'h05c7: oData <= 16'h0000;
            14'h05c8: oData <= 16'h0000;
            14'h05c9: oData <= 16'h0000;
            14'h05ca: oData <= 16'h0000;
            14'h05cb: oData <= 16'h0000;
            14'h05cc: oData <= 16'h0000;
            14'h05cd: oData <= 16'h0aa8;
            14'h05ce: oData <= 16'h0000;
            14'h05cf: oData <= 16'h0000;
            14'h05d0: oData <= 16'h0000;
            14'h05d1: oData <= 16'ha2aa;
            14'h05d2: oData <= 16'haaaa;
            14'h05d3: oData <= 16'hffff;
            14'h05d4: oData <= 16'hffff;
            14'h05d5: oData <= 16'hffff;
            14'h05d6: oData <= 16'haaff;
            14'h05d7: oData <= 16'h0000;
            14'h05d8: oData <= 16'h02aa;
            14'h05d9: oData <= 16'h0000;
            14'h05da: oData <= 16'h0000;
            14'h05db: oData <= 16'h0000;
            14'h05dc: oData <= 16'h0000;
            14'h05dd: oData <= 16'h0000;
            14'h05de: oData <= 16'h0000;
            14'h05df: oData <= 16'h0000;
            14'h05e0: oData <= 16'h0000;
            14'h05e1: oData <= 16'h2aa8;
            14'h05e2: oData <= 16'h0000;
            14'h05e3: oData <= 16'h0000;
            14'h05e4: oData <= 16'h0000;
            14'h05e5: oData <= 16'h02aa;
            14'h05e6: oData <= 16'haa80;
            14'h05e7: oData <= 16'hffaa;
            14'h05e8: oData <= 16'hffff;
            14'h05e9: oData <= 16'hffff;
            14'h05ea: oData <= 16'h2abf;
            14'h05eb: oData <= 16'h8000;
            14'h05ec: oData <= 16'h02aa;
            14'h05ed: oData <= 16'h0000;
            14'h05ee: oData <= 16'h0000;
            14'h05ef: oData <= 16'h0000;
            14'h05f0: oData <= 16'h0000;
            14'h05f1: oData <= 16'h0000;
            14'h05f2: oData <= 16'h0000;
            14'h05f3: oData <= 16'h0000;
            14'h05f4: oData <= 16'h0000;
            14'h05f5: oData <= 16'haaa0;
            14'h05f6: oData <= 16'h0000;
            14'h05f7: oData <= 16'h0000;
            14'h05f8: oData <= 16'h8000;
            14'h05f9: oData <= 16'h02aa;
            14'h05fa: oData <= 16'h8000;
            14'h05fb: oData <= 16'haaaa;
            14'h05fc: oData <= 16'hffff;
            14'h05fd: oData <= 16'hffff;
            14'h05fe: oData <= 16'h02aa;
            14'h05ff: oData <= 16'h8000;
            14'h0600: oData <= 16'h00aa;
            14'h0601: oData <= 16'h0000;
            14'h0602: oData <= 16'h0000;
            14'h0603: oData <= 16'h0000;
            14'h0604: oData <= 16'h0000;
            14'h0605: oData <= 16'h0000;
            14'h0606: oData <= 16'h0000;
            14'h0607: oData <= 16'h0000;
            14'h0608: oData <= 16'h0000;
            14'h0609: oData <= 16'haa80;
            14'h060a: oData <= 16'h0002;
            14'h060b: oData <= 16'h0000;
            14'h060c: oData <= 16'h8000;
            14'h060d: oData <= 16'h00aa;
            14'h060e: oData <= 16'h0000;
            14'h060f: oData <= 16'haa80;
            14'h0610: oData <= 16'haaaa;
            14'h0611: oData <= 16'haaaa;
            14'h0612: oData <= 16'h002a;
            14'h0613: oData <= 16'ha000;
            14'h0614: oData <= 16'h002a;
            14'h0615: oData <= 16'h0000;
            14'h0616: oData <= 16'h0000;
            14'h0617: oData <= 16'h0000;
            14'h0618: oData <= 16'h0000;
            14'h0619: oData <= 16'h0000;
            14'h061a: oData <= 16'h0000;
            14'h061b: oData <= 16'h0000;
            14'h061c: oData <= 16'h0000;
            14'h061d: oData <= 16'haa00;
            14'h061e: oData <= 16'h000a;
            14'h061f: oData <= 16'h0000;
            14'h0620: oData <= 16'h8000;
            14'h0621: oData <= 16'h00aa;
            14'h0622: oData <= 16'h0000;
            14'h0623: oData <= 16'h8000;
            14'h0624: oData <= 16'haaaa;
            14'h0625: oData <= 16'haaaa;
            14'h0626: oData <= 16'h0002;
            14'h0627: oData <= 16'ha800;
            14'h0628: oData <= 16'h002a;
            14'h0629: oData <= 16'h0000;
            14'h062a: oData <= 16'h0000;
            14'h062b: oData <= 16'h0000;
            14'h062c: oData <= 16'h0000;
            14'h062d: oData <= 16'h0000;
            14'h062e: oData <= 16'h0000;
            14'h062f: oData <= 16'h0000;
            14'h0630: oData <= 16'h0000;
            14'h0631: oData <= 16'ha800;
            14'h0632: oData <= 16'h000a;
            14'h0633: oData <= 16'h0000;
            14'h0634: oData <= 16'h8000;
            14'h0635: oData <= 16'h00aa;
            14'h0636: oData <= 16'h0000;
            14'h0637: oData <= 16'h0000;
            14'h0638: oData <= 16'h0000;
            14'h0639: oData <= 16'h0000;
            14'h063a: oData <= 16'h0000;
            14'h063b: oData <= 16'haa00;
            14'h063c: oData <= 16'h000a;
            14'h063d: oData <= 16'h0000;
            14'h063e: oData <= 16'h0000;
            14'h063f: oData <= 16'h0000;
            14'h0640: oData <= 16'h0000;
            14'h0641: oData <= 16'h0000;
            14'h0642: oData <= 16'h0000;
            14'h0643: oData <= 16'h0000;
            14'h0644: oData <= 16'h0000;
            14'h0645: oData <= 16'ha800;
            14'h0646: oData <= 16'h002a;
            14'h0647: oData <= 16'h0000;
            14'h0648: oData <= 16'ha000;
            14'h0649: oData <= 16'h00aa;
            14'h064a: oData <= 16'h0000;
            14'h064b: oData <= 16'h0000;
            14'h064c: oData <= 16'h0000;
            14'h064d: oData <= 16'h0000;
            14'h064e: oData <= 16'h0000;
            14'h064f: oData <= 16'haaa0;
            14'h0650: oData <= 16'h0002;
            14'h0651: oData <= 16'h0000;
            14'h0652: oData <= 16'h0000;
            14'h0653: oData <= 16'h0000;
            14'h0654: oData <= 16'h0000;
            14'h0655: oData <= 16'h0000;
            14'h0656: oData <= 16'h0000;
            14'h0657: oData <= 16'h0000;
            14'h0658: oData <= 16'h0000;
            14'h0659: oData <= 16'ha000;
            14'h065a: oData <= 16'h00aa;
            14'h065b: oData <= 16'h0000;
            14'h065c: oData <= 16'ha000;
            14'h065d: oData <= 16'h002a;
            14'h065e: oData <= 16'h0000;
            14'h065f: oData <= 16'h0000;
            14'h0660: oData <= 16'h0000;
            14'h0661: oData <= 16'h0000;
            14'h0662: oData <= 16'h0000;
            14'h0663: oData <= 16'haaa8;
            14'h0664: oData <= 16'h0002;
            14'h0665: oData <= 16'h0000;
            14'h0666: oData <= 16'h0000;
            14'h0667: oData <= 16'h0000;
            14'h0668: oData <= 16'h0000;
            14'h0669: oData <= 16'h0000;
            14'h066a: oData <= 16'h0000;
            14'h066b: oData <= 16'h0000;
            14'h066c: oData <= 16'h0000;
            14'h066d: oData <= 16'h8000;
            14'h066e: oData <= 16'haaaa;
            14'h066f: oData <= 16'h000a;
            14'h0670: oData <= 16'ha000;
            14'h0671: oData <= 16'h002a;
            14'h0672: oData <= 16'h0000;
            14'h0673: oData <= 16'ha000;
            14'h0674: oData <= 16'h0002;
            14'h0675: oData <= 16'h0000;
            14'h0676: oData <= 16'h0000;
            14'h0677: oData <= 16'h2aa8;
            14'h0678: oData <= 16'h0000;
            14'h0679: oData <= 16'h0000;
            14'h067a: oData <= 16'h0000;
            14'h067b: oData <= 16'h0000;
            14'h067c: oData <= 16'h0000;
            14'h067d: oData <= 16'h0000;
            14'h067e: oData <= 16'h0000;
            14'h067f: oData <= 16'h0000;
            14'h0680: oData <= 16'h0000;
            14'h0681: oData <= 16'h0000;
            14'h0682: oData <= 16'haaaa;
            14'h0683: oData <= 16'haaaa;
            14'h0684: oData <= 16'ha000;
            14'h0685: oData <= 16'h002a;
            14'h0686: oData <= 16'haa80;
            14'h0687: oData <= 16'haaaa;
            14'h0688: oData <= 16'h000a;
            14'h0689: oData <= 16'h0000;
            14'h068a: oData <= 16'h0000;
            14'h068b: oData <= 16'h0aa8;
            14'h068c: oData <= 16'h0000;
            14'h068d: oData <= 16'h0000;
            14'h068e: oData <= 16'h0000;
            14'h068f: oData <= 16'h0000;
            14'h0690: oData <= 16'h0000;
            14'h0691: oData <= 16'h0000;
            14'h0692: oData <= 16'h0000;
            14'h0693: oData <= 16'h0000;
            14'h0694: oData <= 16'h0000;
            14'h0695: oData <= 16'h0000;
            14'h0696: oData <= 16'haaaa;
            14'h0697: oData <= 16'haaaa;
            14'h0698: oData <= 16'haaaa;
            14'h0699: oData <= 16'haaaa;
            14'h069a: oData <= 16'haaaa;
            14'h069b: oData <= 16'haaaa;
            14'h069c: oData <= 16'h002a;
            14'h069d: oData <= 16'h0000;
            14'h069e: oData <= 16'h0000;
            14'h069f: oData <= 16'h0aa8;
            14'h06a0: oData <= 16'h0000;
            14'h06a1: oData <= 16'h0000;
            14'h06a2: oData <= 16'h0000;
            14'h06a3: oData <= 16'h0000;
            14'h06a4: oData <= 16'h0000;
            14'h06a5: oData <= 16'h0000;
            14'h06a6: oData <= 16'h0000;
            14'h06a7: oData <= 16'h0000;
            14'h06a8: oData <= 16'h0000;
            14'h06a9: oData <= 16'h0000;
            14'h06aa: oData <= 16'haaa8;
            14'h06ab: oData <= 16'haaaa;
            14'h06ac: oData <= 16'haaaa;
            14'h06ad: oData <= 16'haaaa;
            14'h06ae: oData <= 16'haaaa;
            14'h06af: oData <= 16'haaaa;
            14'h06b0: oData <= 16'h02aa;
            14'h06b1: oData <= 16'h0000;
            14'h06b2: oData <= 16'h0000;
            14'h06b3: oData <= 16'h2aa8;
            14'h06b4: oData <= 16'h0000;
            14'h06b5: oData <= 16'h0000;
            14'h06b6: oData <= 16'h0000;
            14'h06b7: oData <= 16'h0000;
            14'h06b8: oData <= 16'h0000;
            14'h06b9: oData <= 16'h0000;
            14'h06ba: oData <= 16'h0000;
            14'h06bb: oData <= 16'h0000;
            14'h06bc: oData <= 16'h0000;
            14'h06bd: oData <= 16'h0000;
            14'h06be: oData <= 16'haaa0;
            14'h06bf: oData <= 16'haaaa;
            14'h06c0: oData <= 16'haaaa;
            14'h06c1: oData <= 16'haaaa;
            14'h06c2: oData <= 16'haaaa;
            14'h06c3: oData <= 16'haaaa;
            14'h06c4: oData <= 16'h0aaa;
            14'h06c5: oData <= 16'h0000;
            14'h06c6: oData <= 16'h0000;
            14'h06c7: oData <= 16'haaa0;
            14'h06c8: oData <= 16'h0000;
            14'h06c9: oData <= 16'ha000;
            14'h06ca: oData <= 16'h00aa;
            14'h06cb: oData <= 16'h0000;
            14'h06cc: oData <= 16'h0000;
            14'h06cd: oData <= 16'h0000;
            14'h06ce: oData <= 16'h0000;
            14'h06cf: oData <= 16'h0000;
            14'h06d0: oData <= 16'h0000;
            14'h06d1: oData <= 16'h0000;
            14'h06d2: oData <= 16'h0000;
            14'h06d3: oData <= 16'haaa8;
            14'h06d4: oData <= 16'haaaa;
            14'h06d5: oData <= 16'haaaa;
            14'h06d6: oData <= 16'haaaa;
            14'h06d7: oData <= 16'haaaa;
            14'h06d8: oData <= 16'h2aaa;
            14'h06d9: oData <= 16'h0000;
            14'h06da: oData <= 16'h0000;
            14'h06db: oData <= 16'haa80;
            14'h06dc: oData <= 16'h0002;
            14'h06dd: oData <= 16'haa80;
            14'h06de: oData <= 16'h02aa;
            14'h06df: oData <= 16'h0000;
            14'h06e0: oData <= 16'h0000;
            14'h06e1: oData <= 16'h0000;
            14'h06e2: oData <= 16'h0000;
            14'h06e3: oData <= 16'h0000;
            14'h06e4: oData <= 16'h0000;
            14'h06e5: oData <= 16'h0000;
            14'h06e6: oData <= 16'h0000;
            14'h06e7: oData <= 16'h8000;
            14'h06e8: oData <= 16'haaaa;
            14'h06e9: oData <= 16'haaaa;
            14'h06ea: oData <= 16'h00aa;
            14'h06eb: oData <= 16'h0000;
            14'h06ec: oData <= 16'haaa8;
            14'h06ed: oData <= 16'h0002;
            14'h06ee: oData <= 16'h0000;
            14'h06ef: oData <= 16'haa00;
            14'h06f0: oData <= 16'h000a;
            14'h06f1: oData <= 16'haaa0;
            14'h06f2: oData <= 16'h0aaa;
            14'h06f3: oData <= 16'h0000;
            14'h06f4: oData <= 16'h0000;
            14'h06f5: oData <= 16'h0000;
            14'h06f6: oData <= 16'h0000;
            14'h06f7: oData <= 16'h0000;
            14'h06f8: oData <= 16'h0000;
            14'h06f9: oData <= 16'h0000;
            14'h06fa: oData <= 16'h0000;
            14'h06fb: oData <= 16'h0000;
            14'h06fc: oData <= 16'haa00;
            14'h06fd: oData <= 16'h0002;
            14'h06fe: oData <= 16'h0000;
            14'h06ff: oData <= 16'h0000;
            14'h0700: oData <= 16'haaa0;
            14'h0701: oData <= 16'h000a;
            14'h0702: oData <= 16'h0000;
            14'h0703: oData <= 16'ha800;
            14'h0704: oData <= 16'h002a;
            14'h0705: oData <= 16'haaa8;
            14'h0706: oData <= 16'h2aaa;
            14'h0707: oData <= 16'h0000;
            14'h0708: oData <= 16'h0000;
            14'h0709: oData <= 16'h0000;
            14'h070a: oData <= 16'h0000;
            14'h070b: oData <= 16'h0000;
            14'h070c: oData <= 16'h0000;
            14'h070d: oData <= 16'h0000;
            14'h070e: oData <= 16'h0000;
            14'h070f: oData <= 16'h0000;
            14'h0710: oData <= 16'haa00;
            14'h0711: oData <= 16'h0002;
            14'h0712: oData <= 16'h0000;
            14'h0713: oData <= 16'h0000;
            14'h0714: oData <= 16'haa00;
            14'h0715: oData <= 16'h002a;
            14'h0716: oData <= 16'h0000;
            14'h0717: oData <= 16'ha000;
            14'h0718: oData <= 16'h00aa;
            14'h0719: oData <= 16'h2aa8;
            14'h071a: oData <= 16'h2aa0;
            14'h071b: oData <= 16'h0000;
            14'h071c: oData <= 16'h0000;
            14'h071d: oData <= 16'h0000;
            14'h071e: oData <= 16'h0000;
            14'h071f: oData <= 16'h0000;
            14'h0720: oData <= 16'h0000;
            14'h0721: oData <= 16'h0000;
            14'h0722: oData <= 16'h0000;
            14'h0723: oData <= 16'h0000;
            14'h0724: oData <= 16'haa00;
            14'h0725: oData <= 16'h0002;
            14'h0726: oData <= 16'h0000;
            14'h0727: oData <= 16'h0000;
            14'h0728: oData <= 16'ha800;
            14'h0729: oData <= 16'h02aa;
            14'h072a: oData <= 16'h0000;
            14'h072b: oData <= 16'h8000;
            14'h072c: oData <= 16'h00aa;
            14'h072d: oData <= 16'h02aa;
            14'h072e: oData <= 16'h2aa0;
            14'h072f: oData <= 16'h0000;
            14'h0730: oData <= 16'h0000;
            14'h0731: oData <= 16'h0000;
            14'h0732: oData <= 16'h0000;
            14'h0733: oData <= 16'h0000;
            14'h0734: oData <= 16'h0000;
            14'h0735: oData <= 16'h0000;
            14'h0736: oData <= 16'h0000;
            14'h0737: oData <= 16'h0000;
            14'h0738: oData <= 16'haa80;
            14'h0739: oData <= 16'h0002;
            14'h073a: oData <= 16'h0000;
            14'h073b: oData <= 16'h0000;
            14'h073c: oData <= 16'ha000;
            14'h073d: oData <= 16'h0aaa;
            14'h073e: oData <= 16'h0000;
            14'h073f: oData <= 16'h0000;
            14'h0740: oData <= 16'h00aa;
            14'h0741: oData <= 16'h02aa;
            14'h0742: oData <= 16'h2aa0;
            14'h0743: oData <= 16'h0000;
            14'h0744: oData <= 16'h0000;
            14'h0745: oData <= 16'h0000;
            14'h0746: oData <= 16'h0000;
            14'h0747: oData <= 16'h0000;
            14'h0748: oData <= 16'h0000;
            14'h0749: oData <= 16'h0000;
            14'h074a: oData <= 16'h0000;
            14'h074b: oData <= 16'h0000;
            14'h074c: oData <= 16'haa80;
            14'h074d: oData <= 16'h0000;
            14'h074e: oData <= 16'h0000;
            14'h074f: oData <= 16'h0000;
            14'h0750: oData <= 16'h0000;
            14'h0751: oData <= 16'haaaa;
            14'h0752: oData <= 16'h0000;
            14'h0753: oData <= 16'h0000;
            14'h0754: oData <= 16'h0028;
            14'h0755: oData <= 16'h00aa;
            14'h0756: oData <= 16'h0aa8;
            14'h0757: oData <= 16'h0000;
            14'h0758: oData <= 16'h0000;
            14'h0759: oData <= 16'h0000;
            14'h075a: oData <= 16'h0000;
            14'h075b: oData <= 16'h0000;
            14'h075c: oData <= 16'h0000;
            14'h075d: oData <= 16'h0000;
            14'h075e: oData <= 16'h0000;
            14'h075f: oData <= 16'h0000;
            14'h0760: oData <= 16'haa80;
            14'h0761: oData <= 16'h0000;
            14'h0762: oData <= 16'h0000;
            14'h0763: oData <= 16'h0000;
            14'h0764: oData <= 16'h0000;
            14'h0765: oData <= 16'haaa8;
            14'h0766: oData <= 16'h0002;
            14'h0767: oData <= 16'h0000;
            14'h0768: oData <= 16'h0000;
            14'h0769: oData <= 16'h00aa;
            14'h076a: oData <= 16'h0aa8;
            14'h076b: oData <= 16'h0280;
            14'h076c: oData <= 16'h0000;
            14'h076d: oData <= 16'h0000;
            14'h076e: oData <= 16'h0000;
            14'h076f: oData <= 16'h0000;
            14'h0770: oData <= 16'h0000;
            14'h0771: oData <= 16'h0000;
            14'h0772: oData <= 16'h0000;
            14'h0773: oData <= 16'h0000;
            14'h0774: oData <= 16'haa80;
            14'h0775: oData <= 16'h0000;
            14'h0776: oData <= 16'h0000;
            14'h0777: oData <= 16'h0000;
            14'h0778: oData <= 16'h0000;
            14'h0779: oData <= 16'haaa0;
            14'h077a: oData <= 16'h0002;
            14'h077b: oData <= 16'h0000;
            14'h077c: oData <= 16'h0000;
            14'h077d: oData <= 16'ha0aa;
            14'h077e: oData <= 16'h02aa;
            14'h077f: oData <= 16'h0aa0;
            14'h0780: oData <= 16'h0000;
            14'h0781: oData <= 16'h0000;
            14'h0782: oData <= 16'h0000;
            14'h0783: oData <= 16'h0000;
            14'h0784: oData <= 16'h0000;
            14'h0785: oData <= 16'h0000;
            14'h0786: oData <= 16'h0000;
            14'h0787: oData <= 16'h0000;
            14'h0788: oData <= 16'haaa0;
            14'h0789: oData <= 16'h0000;
            14'h078a: oData <= 16'h0000;
            14'h078b: oData <= 16'h0000;
            14'h078c: oData <= 16'h0000;
            14'h078d: oData <= 16'haa00;
            14'h078e: oData <= 16'h0002;
            14'h078f: oData <= 16'h0000;
            14'h0790: oData <= 16'h0000;
            14'h0791: oData <= 16'haaaa;
            14'h0792: oData <= 16'h02aa;
            14'h0793: oData <= 16'h0aa0;
            14'h0794: oData <= 16'h0000;
            14'h0795: oData <= 16'h0000;
            14'h0796: oData <= 16'h0000;
            14'h0797: oData <= 16'h0000;
            14'h0798: oData <= 16'h0000;
            14'h0799: oData <= 16'h0000;
            14'h079a: oData <= 16'h0000;
            14'h079b: oData <= 16'h0000;
            14'h079c: oData <= 16'h2aa0;
            14'h079d: oData <= 16'h0000;
            14'h079e: oData <= 16'h0000;
            14'h079f: oData <= 16'h0000;
            14'h07a0: oData <= 16'h0000;
            14'h07a1: oData <= 16'ha800;
            14'h07a2: oData <= 16'h0000;
            14'h07a3: oData <= 16'h0000;
            14'h07a4: oData <= 16'h0000;
            14'h07a5: oData <= 16'haaaa;
            14'h07a6: oData <= 16'h00aa;
            14'h07a7: oData <= 16'h0aa8;
            14'h07a8: oData <= 16'h0000;
            14'h07a9: oData <= 16'h0000;
            14'h07aa: oData <= 16'h0000;
            14'h07ab: oData <= 16'h00a8;
            14'h07ac: oData <= 16'h0000;
            14'h07ad: oData <= 16'h0000;
            14'h07ae: oData <= 16'h0000;
            14'h07af: oData <= 16'h0000;
            14'h07b0: oData <= 16'h2aa0;
            14'h07b1: oData <= 16'h0000;
            14'h07b2: oData <= 16'h0000;
            14'h07b3: oData <= 16'h0000;
            14'h07b4: oData <= 16'h0000;
            14'h07b5: oData <= 16'h0000;
            14'h07b6: oData <= 16'h0000;
            14'h07b7: oData <= 16'h0000;
            14'h07b8: oData <= 16'h0000;
            14'h07b9: oData <= 16'haaa8;
            14'h07ba: oData <= 16'h000a;
            14'h07bb: oData <= 16'h0aa8;
            14'h07bc: oData <= 16'h0000;
            14'h07bd: oData <= 16'h0000;
            14'h07be: oData <= 16'h0000;
            14'h07bf: oData <= 16'h02aa;
            14'h07c0: oData <= 16'h0000;
            14'h07c1: oData <= 16'h0000;
            14'h07c2: oData <= 16'h0000;
            14'h07c3: oData <= 16'h0000;
            14'h07c4: oData <= 16'h2aa0;
            14'h07c5: oData <= 16'h0000;
            14'h07c6: oData <= 16'h0000;
            14'h07c7: oData <= 16'h0000;
            14'h07c8: oData <= 16'h0000;
            14'h07c9: oData <= 16'h0000;
            14'h07ca: oData <= 16'h0000;
            14'h07cb: oData <= 16'h0000;
            14'h07cc: oData <= 16'h0000;
            14'h07cd: oData <= 16'haaa0;
            14'h07ce: oData <= 16'h0000;
            14'h07cf: oData <= 16'h02aa;
            14'h07d0: oData <= 16'h0000;
            14'h07d1: oData <= 16'h0000;
            14'h07d2: oData <= 16'h0000;
            14'h07d3: oData <= 16'h2aaa;
            14'h07d4: oData <= 16'h0000;
            14'h07d5: oData <= 16'h0000;
            14'h07d6: oData <= 16'h0000;
            14'h07d7: oData <= 16'h0000;
            14'h07d8: oData <= 16'h2aa8;
            14'h07d9: oData <= 16'h0000;
            14'h07da: oData <= 16'h0000;
            14'h07db: oData <= 16'h0000;
            14'h07dc: oData <= 16'h0000;
            14'h07dd: oData <= 16'h0000;
            14'h07de: oData <= 16'h0000;
            14'h07df: oData <= 16'h0000;
            14'h07e0: oData <= 16'h0000;
            14'h07e1: oData <= 16'h0000;
            14'h07e2: oData <= 16'h8000;
            14'h07e3: oData <= 16'h02aa;
            14'h07e4: oData <= 16'h0000;
            14'h07e5: oData <= 16'h0000;
            14'h07e6: oData <= 16'h0000;
            14'h07e7: oData <= 16'haaaa;
            14'h07e8: oData <= 16'h0002;
            14'h07e9: oData <= 16'h0000;
            14'h07ea: oData <= 16'h0000;
            14'h07eb: oData <= 16'h0000;
            14'h07ec: oData <= 16'h0aa8;
            14'h07ed: oData <= 16'h0000;
            14'h07ee: oData <= 16'h0000;
            14'h07ef: oData <= 16'h0000;
            14'h07f0: oData <= 16'h0000;
            14'h07f1: oData <= 16'h0000;
            14'h07f2: oData <= 16'h0000;
            14'h07f3: oData <= 16'h0000;
            14'h07f4: oData <= 16'h0000;
            14'h07f5: oData <= 16'h0000;
            14'h07f6: oData <= 16'ha000;
            14'h07f7: oData <= 16'h00aa;
            14'h07f8: oData <= 16'h0000;
            14'h07f9: oData <= 16'h0000;
            14'h07fa: oData <= 16'h0000;
            14'h07fb: oData <= 16'haaa8;
            14'h07fc: oData <= 16'h000a;
            14'h07fd: oData <= 16'h0000;
            14'h07fe: oData <= 16'h0000;
            14'h07ff: oData <= 16'h0000;
            14'h0800: oData <= 16'h0aaa;
            14'h0801: oData <= 16'h0000;
            14'h0802: oData <= 16'h0000;
            14'h0803: oData <= 16'h0000;
            14'h0804: oData <= 16'h0000;
            14'h0805: oData <= 16'h0000;
            14'h0806: oData <= 16'h0000;
            14'h0807: oData <= 16'h0000;
            14'h0808: oData <= 16'h0000;
            14'h0809: oData <= 16'h0000;
            14'h080a: oData <= 16'haa80;
            14'h080b: oData <= 16'h002a;
            14'h080c: oData <= 16'h0000;
            14'h080d: oData <= 16'h0000;
            14'h080e: oData <= 16'h0000;
            14'h080f: oData <= 16'haaa0;
            14'h0810: oData <= 16'h00aa;
            14'h0811: oData <= 16'h0000;
            14'h0812: oData <= 16'h0000;
            14'h0813: oData <= 16'h8000;
            14'h0814: oData <= 16'h0aaa;
            14'h0815: oData <= 16'h0000;
            14'h0816: oData <= 16'h0000;
            14'h0817: oData <= 16'h0000;
            14'h0818: oData <= 16'h0000;
            14'h0819: oData <= 16'h0000;
            14'h081a: oData <= 16'h0000;
            14'h081b: oData <= 16'h0000;
            14'h081c: oData <= 16'h0000;
            14'h081d: oData <= 16'h0000;
            14'h081e: oData <= 16'haaaa;
            14'h081f: oData <= 16'h000a;
            14'h0820: oData <= 16'h0000;
            14'h0821: oData <= 16'h0000;
            14'h0822: oData <= 16'h0000;
            14'h0823: oData <= 16'haa00;
            14'h0824: oData <= 16'h0aaa;
            14'h0825: oData <= 16'h0000;
            14'h0826: oData <= 16'h0000;
            14'h0827: oData <= 16'haa80;
            14'h0828: oData <= 16'haaaa;
            14'h0829: oData <= 16'haaaa;
            14'h082a: oData <= 16'haaaa;
            14'h082b: oData <= 16'h0aaa;
            14'h082c: oData <= 16'h0000;
            14'h082d: oData <= 16'h0000;
            14'h082e: oData <= 16'h0000;
            14'h082f: oData <= 16'h0000;
            14'h0830: oData <= 16'h0000;
            14'h0831: oData <= 16'h8000;
            14'h0832: oData <= 16'haaaa;
            14'h0833: oData <= 16'h0002;
            14'h0834: oData <= 16'h0000;
            14'h0835: oData <= 16'h0000;
            14'h0836: oData <= 16'h0000;
            14'h0837: oData <= 16'ha000;
            14'h0838: oData <= 16'h2aaa;
            14'h0839: oData <= 16'h0000;
            14'h083a: oData <= 16'h8000;
            14'h083b: oData <= 16'haaaa;
            14'h083c: oData <= 16'haaaa;
            14'h083d: oData <= 16'haaaa;
            14'h083e: oData <= 16'haaaa;
            14'h083f: oData <= 16'h2aaa;
            14'h0840: oData <= 16'h0000;
            14'h0841: oData <= 16'h0000;
            14'h0842: oData <= 16'h0000;
            14'h0843: oData <= 16'h0000;
            14'h0844: oData <= 16'h0000;
            14'h0845: oData <= 16'h8000;
            14'h0846: oData <= 16'h2aaa;
            14'h0847: oData <= 16'h0000;
            14'h0848: oData <= 16'h0000;
            14'h0849: oData <= 16'h0000;
            14'h084a: oData <= 16'h0000;
            14'h084b: oData <= 16'h0000;
            14'h084c: oData <= 16'haaaa;
            14'h084d: oData <= 16'h0002;
            14'h084e: oData <= 16'haa80;
            14'h084f: oData <= 16'haaaa;
            14'h0850: oData <= 16'haaaa;
            14'h0851: oData <= 16'haaaa;
            14'h0852: oData <= 16'haaaa;
            14'h0853: oData <= 16'haaaa;
            14'h0854: oData <= 16'h0000;
            14'h0855: oData <= 16'h0000;
            14'h0856: oData <= 16'h0000;
            14'h0857: oData <= 16'h0000;
            14'h0858: oData <= 16'h0000;
            14'h0859: oData <= 16'ha000;
            14'h085a: oData <= 16'h02aa;
            14'h085b: oData <= 16'h0000;
            14'h085c: oData <= 16'h0000;
            14'h085d: oData <= 16'h0000;
            14'h085e: oData <= 16'h0000;
            14'h085f: oData <= 16'h0000;
            14'h0860: oData <= 16'haaa8;
            14'h0861: oData <= 16'h802a;
            14'h0862: oData <= 16'haaaa;
            14'h0863: oData <= 16'haaaa;
            14'h0864: oData <= 16'haaaa;
            14'h0865: oData <= 16'haaaa;
            14'h0866: oData <= 16'haaaa;
            14'h0867: oData <= 16'haaaa;
            14'h0868: oData <= 16'h000a;
            14'h0869: oData <= 16'h0000;
            14'h086a: oData <= 16'h0000;
            14'h086b: oData <= 16'h0000;
            14'h086c: oData <= 16'h0000;
            14'h086d: oData <= 16'ha000;
            14'h086e: oData <= 16'h002a;
            14'h086f: oData <= 16'h0000;
            14'h0870: oData <= 16'h0000;
            14'h0871: oData <= 16'h0000;
            14'h0872: oData <= 16'h0000;
            14'h0873: oData <= 16'h0000;
            14'h0874: oData <= 16'haa80;
            14'h0875: oData <= 16'haaaa;
            14'h0876: oData <= 16'haaaa;
            14'h0877: oData <= 16'haaaa;
            14'h0878: oData <= 16'haaaa;
            14'h0879: oData <= 16'haaaa;
            14'h087a: oData <= 16'haaaa;
            14'h087b: oData <= 16'haaaa;
            14'h087c: oData <= 16'h002a;
            14'h087d: oData <= 16'h0000;
            14'h087e: oData <= 16'h0000;
            14'h087f: oData <= 16'h0000;
            14'h0880: oData <= 16'h0000;
            14'h0881: oData <= 16'ha000;
            14'h0882: oData <= 16'h002a;
            14'h0883: oData <= 16'h0000;
            14'h0884: oData <= 16'h0000;
            14'h0885: oData <= 16'h0000;
            14'h0886: oData <= 16'h0000;
            14'h0887: oData <= 16'h0000;
            14'h0888: oData <= 16'ha800;
            14'h0889: oData <= 16'haaaa;
            14'h088a: oData <= 16'haaaa;
            14'h088b: oData <= 16'h00aa;
            14'h088c: oData <= 16'h0000;
            14'h088d: oData <= 16'h0000;
            14'h088e: oData <= 16'h0000;
            14'h088f: oData <= 16'haa00;
            14'h0890: oData <= 16'h00aa;
            14'h0891: oData <= 16'h0000;
            14'h0892: oData <= 16'h0000;
            14'h0893: oData <= 16'h0000;
            14'h0894: oData <= 16'h0000;
            14'h0895: oData <= 16'ha000;
            14'h0896: oData <= 16'h002a;
            14'h0897: oData <= 16'h0000;
            14'h0898: oData <= 16'h0000;
            14'h0899: oData <= 16'h0000;
            14'h089a: oData <= 16'h0000;
            14'h089b: oData <= 16'h0000;
            14'h089c: oData <= 16'ha000;
            14'h089d: oData <= 16'haaaa;
            14'h089e: oData <= 16'haaaa;
            14'h089f: oData <= 16'h0000;
            14'h08a0: oData <= 16'h0000;
            14'h08a1: oData <= 16'h0000;
            14'h08a2: oData <= 16'h0000;
            14'h08a3: oData <= 16'ha000;
            14'h08a4: oData <= 16'h0aaa;
            14'h08a5: oData <= 16'h0000;
            14'h08a6: oData <= 16'h0000;
            14'h08a7: oData <= 16'h0000;
            14'h08a8: oData <= 16'h0000;
            14'h08a9: oData <= 16'h8000;
            14'h08aa: oData <= 16'h00aa;
            14'h08ab: oData <= 16'h0000;
            14'h08ac: oData <= 16'h0000;
            14'h08ad: oData <= 16'h0000;
            14'h08ae: oData <= 16'h0000;
            14'h08af: oData <= 16'h0000;
            14'h08b0: oData <= 16'h0000;
            14'h08b1: oData <= 16'haaaa;
            14'h08b2: oData <= 16'h00aa;
            14'h08b3: oData <= 16'h0000;
            14'h08b4: oData <= 16'h0000;
            14'h08b5: oData <= 16'h0000;
            14'h08b6: oData <= 16'h0000;
            14'h08b7: oData <= 16'h8000;
            14'h08b8: oData <= 16'h2aaa;
            14'h08b9: oData <= 16'h0000;
            14'h08ba: oData <= 16'h0000;
            14'h08bb: oData <= 16'h0000;
            14'h08bc: oData <= 16'h0000;
            14'h08bd: oData <= 16'h8000;
            14'h08be: oData <= 16'h02aa;
            14'h08bf: oData <= 16'h0000;
            14'h08c0: oData <= 16'h0000;
            14'h08c1: oData <= 16'h0000;
            14'h08c2: oData <= 16'h0000;
            14'h08c3: oData <= 16'h0000;
            14'h08c4: oData <= 16'h0000;
            14'h08c5: oData <= 16'haaa0;
            14'h08c6: oData <= 16'h0000;
            14'h08c7: oData <= 16'h0000;
            14'h08c8: oData <= 16'h0000;
            14'h08c9: oData <= 16'h0000;
            14'h08ca: oData <= 16'h0000;
            14'h08cb: oData <= 16'h0000;
            14'h08cc: oData <= 16'haaa8;
            14'h08cd: oData <= 16'h0002;
            14'h08ce: oData <= 16'h0000;
            14'h08cf: oData <= 16'h0000;
            14'h08d0: oData <= 16'h0000;
            14'h08d1: oData <= 16'h0000;
            14'h08d2: oData <= 16'h02aa;
            14'h08d3: oData <= 16'h0000;
            14'h08d4: oData <= 16'h0000;
            14'h08d5: oData <= 16'h0000;
            14'h08d6: oData <= 16'h0000;
            14'h08d7: oData <= 16'h0000;
            14'h08d8: oData <= 16'h0000;
            14'h08d9: oData <= 16'h0000;
            14'h08da: oData <= 16'h0000;
            14'h08db: oData <= 16'h0000;
            14'h08dc: oData <= 16'h0000;
            14'h08dd: oData <= 16'h0000;
            14'h08de: oData <= 16'h0000;
            14'h08df: oData <= 16'h0000;
            14'h08e0: oData <= 16'haaa0;
            14'h08e1: oData <= 16'h000a;
            14'h08e2: oData <= 16'h0000;
            14'h08e3: oData <= 16'h0000;
            14'h08e4: oData <= 16'h0000;
            14'h08e5: oData <= 16'h0000;
            14'h08e6: oData <= 16'h0aa8;
            14'h08e7: oData <= 16'h0000;
            14'h08e8: oData <= 16'h0000;
            14'h08e9: oData <= 16'h0000;
            14'h08ea: oData <= 16'h0000;
            14'h08eb: oData <= 16'h0000;
            14'h08ec: oData <= 16'h0000;
            14'h08ed: oData <= 16'h0000;
            14'h08ee: oData <= 16'h0000;
            14'h08ef: oData <= 16'h0000;
            14'h08f0: oData <= 16'h0000;
            14'h08f1: oData <= 16'h0000;
            14'h08f2: oData <= 16'h0000;
            14'h08f3: oData <= 16'h0000;
            14'h08f4: oData <= 16'haa80;
            14'h08f5: oData <= 16'h00aa;
            14'h08f6: oData <= 16'h0000;
            14'h08f7: oData <= 16'h0000;
            14'h08f8: oData <= 16'h0000;
            14'h08f9: oData <= 16'h0000;
            14'h08fa: oData <= 16'h2aa8;
            14'h08fb: oData <= 16'h0000;
            14'h08fc: oData <= 16'h0000;
            14'h08fd: oData <= 16'h0000;
            14'h08fe: oData <= 16'h0000;
            14'h08ff: oData <= 16'h0000;
            14'h0900: oData <= 16'h0000;
            14'h0901: oData <= 16'h0000;
            14'h0902: oData <= 16'h0000;
            14'h0903: oData <= 16'h0000;
            14'h0904: oData <= 16'h0000;
            14'h0905: oData <= 16'h0000;
            14'h0906: oData <= 16'h0000;
            14'h0907: oData <= 16'h0000;
            14'h0908: oData <= 16'ha800;
            14'h0909: oData <= 16'h02aa;
            14'h090a: oData <= 16'h0000;
            14'h090b: oData <= 16'h0000;
            14'h090c: oData <= 16'h0000;
            14'h090d: oData <= 16'h0000;
            14'h090e: oData <= 16'h2aa0;
            14'h090f: oData <= 16'h0000;
            14'h0910: oData <= 16'h0000;
            14'h0911: oData <= 16'h0000;
            14'h0912: oData <= 16'h0000;
            14'h0913: oData <= 16'h0000;
            14'h0914: oData <= 16'h0000;
            14'h0915: oData <= 16'h0000;
            14'h0916: oData <= 16'h0000;
            14'h0917: oData <= 16'h0000;
            14'h0918: oData <= 16'h0000;
            14'h0919: oData <= 16'h0000;
            14'h091a: oData <= 16'h0000;
            14'h091b: oData <= 16'h0000;
            14'h091c: oData <= 16'ha000;
            14'h091d: oData <= 16'h02aa;
            14'h091e: oData <= 16'h0000;
            14'h091f: oData <= 16'h0000;
            14'h0920: oData <= 16'h0000;
            14'h0921: oData <= 16'h0000;
            14'h0922: oData <= 16'h0a80;
            14'h0923: oData <= 16'h0000;
            14'h0924: oData <= 16'h0000;
            14'h0925: oData <= 16'h0000;
            14'h0926: oData <= 16'h0000;
            14'h0927: oData <= 16'h0000;
            14'h0928: oData <= 16'h0000;
            14'h0929: oData <= 16'h0000;
            14'h092a: oData <= 16'h0000;
            14'h092b: oData <= 16'h0000;
            14'h092c: oData <= 16'h0000;
            14'h092d: oData <= 16'h0000;
            14'h092e: oData <= 16'h0000;
            14'h092f: oData <= 16'h0000;
            14'h0930: oData <= 16'h0000;
            14'h0931: oData <= 16'h02aa;
            14'h0932: oData <= 16'h0000;
            14'h0933: oData <= 16'h0000;
            14'h0934: oData <= 16'h0000;
            14'h0935: oData <= 16'h0000;
            14'h0936: oData <= 16'h0000;
            14'h0937: oData <= 16'h0000;
            14'h0938: oData <= 16'h0000;
            14'h0939: oData <= 16'h0000;
            14'h093a: oData <= 16'h0000;
            14'h093b: oData <= 16'h0000;
            14'h093c: oData <= 16'h0000;
            14'h093d: oData <= 16'h0000;
            14'h093e: oData <= 16'h0000;
            14'h093f: oData <= 16'h0000;
            14'h0940: oData <= 16'h0000;
            14'h0941: oData <= 16'h0000;
            14'h0942: oData <= 16'h0000;
            14'h0943: oData <= 16'h0000;
            14'h0944: oData <= 16'h0000;
            14'h0945: oData <= 16'h00a8;
            14'h0946: oData <= 16'h0000;
            14'h0947: oData <= 16'h0000;
            14'h0948: oData <= 16'h0000;
            14'h0949: oData <= 16'h0000;
            14'h094a: oData <= 16'h0000;
            14'h094b: oData <= 16'h0000;
            14'h094c: oData <= 16'h0000;
            14'h094d: oData <= 16'h0000;
            14'h094e: oData <= 16'h0000;
            14'h094f: oData <= 16'h0000;
            14'h0950: oData <= 16'h0000;
            14'h0951: oData <= 16'h0000;
            14'h0952: oData <= 16'h0000;
            14'h0953: oData <= 16'h0000;
            14'h0954: oData <= 16'h0000;
            14'h0955: oData <= 16'h0000;
            14'h0956: oData <= 16'h0000;
            14'h0957: oData <= 16'h0000;
            14'h0958: oData <= 16'h0000;
            14'h0959: oData <= 16'h0000;
            14'h095a: oData <= 16'h0000;
            14'h095b: oData <= 16'h0000;
            14'h095c: oData <= 16'h0000;
            14'h095d: oData <= 16'h0000;
            14'h095e: oData <= 16'h0000;
            14'h095f: oData <= 16'h0000;
            14'h0960: oData <= 16'h0000;
            14'h0961: oData <= 16'h0000;
            14'h0962: oData <= 16'h0000;
            14'h0963: oData <= 16'ha800;
            14'h0964: oData <= 16'h0000;
            14'h0965: oData <= 16'h0000;
            14'h0966: oData <= 16'h0000;
            14'h0967: oData <= 16'h0000;
            14'h0968: oData <= 16'h0000;
            14'h0969: oData <= 16'h0000;
            14'h096a: oData <= 16'h0000;
            14'h096b: oData <= 16'h0000;
            14'h096c: oData <= 16'h0000;
            14'h096d: oData <= 16'h0000;
            14'h096e: oData <= 16'h0000;
            14'h096f: oData <= 16'h0000;
            14'h0970: oData <= 16'h0000;
            14'h0971: oData <= 16'h0000;
            14'h0972: oData <= 16'h0000;
            14'h0973: oData <= 16'h0000;
            14'h0974: oData <= 16'h0000;
            14'h0975: oData <= 16'h0000;
            14'h0976: oData <= 16'h0000;
            14'h0977: oData <= 16'haa00;
            14'h0978: oData <= 16'h0002;
            14'h0979: oData <= 16'h0000;
            14'h097a: oData <= 16'h0000;
            14'h097b: oData <= 16'haa80;
            14'h097c: oData <= 16'haaaa;
            14'h097d: oData <= 16'haaaa;
            14'h097e: oData <= 16'haaaa;
            14'h097f: oData <= 16'h2aaa;
            14'h0980: oData <= 16'h0000;
            14'h0981: oData <= 16'h0000;
            14'h0982: oData <= 16'h0000;
            14'h0983: oData <= 16'h0000;
            14'h0984: oData <= 16'h0000;
            14'h0985: oData <= 16'h0000;
            14'h0986: oData <= 16'h0000;
            14'h0987: oData <= 16'h0000;
            14'h0988: oData <= 16'h0000;
            14'h0989: oData <= 16'h0000;
            14'h098a: oData <= 16'h0000;
            14'h098b: oData <= 16'haa00;
            14'h098c: oData <= 16'h0002;
            14'h098d: oData <= 16'h0000;
            14'h098e: oData <= 16'h0000;
            14'h098f: oData <= 16'haaa8;
            14'h0990: oData <= 16'haaaa;
            14'h0991: oData <= 16'haaaa;
            14'h0992: oData <= 16'haaaa;
            14'h0993: oData <= 16'haaaa;
            14'h0994: oData <= 16'haaaa;
            14'h0995: oData <= 16'h000a;
            14'h0996: oData <= 16'h0000;
            14'h0997: oData <= 16'h0000;
            14'h0998: oData <= 16'h0000;
            14'h0999: oData <= 16'h0000;
            14'h099a: oData <= 16'h0000;
            14'h099b: oData <= 16'h0000;
            14'h099c: oData <= 16'h0000;
            14'h099d: oData <= 16'h0000;
            14'h099e: oData <= 16'h0000;
            14'h099f: oData <= 16'ha800;
            14'h09a0: oData <= 16'h000a;
            14'h09a1: oData <= 16'h0000;
            14'h09a2: oData <= 16'h8000;
            14'h09a3: oData <= 16'hffaa;
            14'h09a4: oData <= 16'hffff;
            14'h09a5: oData <= 16'hffff;
            14'h09a6: oData <= 16'hffff;
            14'h09a7: oData <= 16'hafff;
            14'h09a8: oData <= 16'haaaa;
            14'h09a9: oData <= 16'h0aaa;
            14'h09aa: oData <= 16'h0000;
            14'h09ab: oData <= 16'h0000;
            14'h09ac: oData <= 16'h0000;
            14'h09ad: oData <= 16'h0000;
            14'h09ae: oData <= 16'h0000;
            14'h09af: oData <= 16'h0000;
            14'h09b0: oData <= 16'h0000;
            14'h09b1: oData <= 16'h0000;
            14'h09b2: oData <= 16'h0aa8;
            14'h09b3: oData <= 16'ha800;
            14'h09b4: oData <= 16'h000a;
            14'h09b5: oData <= 16'h0000;
            14'h09b6: oData <= 16'ha000;
            14'h09b7: oData <= 16'hfffa;
            14'h09b8: oData <= 16'hffff;
            14'h09b9: oData <= 16'haaab;
            14'h09ba: oData <= 16'haaaa;
            14'h09bb: oData <= 16'hfffa;
            14'h09bc: oData <= 16'hffff;
            14'h09bd: oData <= 16'haaab;
            14'h09be: oData <= 16'h002a;
            14'h09bf: oData <= 16'h0000;
            14'h09c0: oData <= 16'h0000;
            14'h09c1: oData <= 16'h0000;
            14'h09c2: oData <= 16'h0000;
            14'h09c3: oData <= 16'h0000;
            14'h09c4: oData <= 16'h0000;
            14'h09c5: oData <= 16'h0000;
            14'h09c6: oData <= 16'haaaa;
            14'h09c7: oData <= 16'ha002;
            14'h09c8: oData <= 16'h002a;
            14'h09c9: oData <= 16'h0000;
            14'h09ca: oData <= 16'ha800;
            14'h09cb: oData <= 16'hffff;
            14'h09cc: oData <= 16'hafff;
            14'h09cd: oData <= 16'hfffe;
            14'h09ce: oData <= 16'hffff;
            14'h09cf: oData <= 16'haaaf;
            14'h09d0: oData <= 16'haaaa;
            14'h09d1: oData <= 16'habfa;
            14'h09d2: oData <= 16'h02aa;
            14'h09d3: oData <= 16'h0000;
            14'h09d4: oData <= 16'h0000;
            14'h09d5: oData <= 16'h0000;
            14'h09d6: oData <= 16'h0000;
            14'h09d7: oData <= 16'h0000;
            14'h09d8: oData <= 16'h0000;
            14'h09d9: oData <= 16'h0000;
            14'h09da: oData <= 16'haaaa;
            14'h09db: oData <= 16'ha00a;
            14'h09dc: oData <= 16'h002a;
            14'h09dd: oData <= 16'h000a;
            14'h09de: oData <= 16'hea00;
            14'h09df: oData <= 16'hffff;
            14'h09e0: oData <= 16'hfaff;
            14'h09e1: oData <= 16'hafff;
            14'h09e2: oData <= 16'hfeaa;
            14'h09e3: oData <= 16'hffff;
            14'h09e4: oData <= 16'hffff;
            14'h09e5: oData <= 16'hffff;
            14'h09e6: oData <= 16'h0aaf;
            14'h09e7: oData <= 16'h0000;
            14'h09e8: oData <= 16'h0000;
            14'h09e9: oData <= 16'h0000;
            14'h09ea: oData <= 16'h0000;
            14'h09eb: oData <= 16'h0000;
            14'h09ec: oData <= 16'h0000;
            14'h09ed: oData <= 16'h8000;
            14'h09ee: oData <= 16'haaaa;
            14'h09ef: oData <= 16'h802a;
            14'h09f0: oData <= 16'ha0aa;
            14'h09f1: oData <= 16'h002a;
            14'h09f2: oData <= 16'hfa00;
            14'h09f3: oData <= 16'hffff;
            14'h09f4: oData <= 16'hffaf;
            14'h09f5: oData <= 16'hfaab;
            14'h09f6: oData <= 16'habff;
            14'h09f7: oData <= 16'hfffe;
            14'h09f8: oData <= 16'hffff;
            14'h09f9: oData <= 16'haaaf;
            14'h09fa: oData <= 16'haaff;
            14'h09fb: oData <= 16'h0000;
            14'h09fc: oData <= 16'h0000;
            14'h09fd: oData <= 16'h0000;
            14'h09fe: oData <= 16'h0000;
            14'h09ff: oData <= 16'h0000;
            14'h0a00: oData <= 16'h0000;
            14'h0a01: oData <= 16'ha000;
            14'h0a02: oData <= 16'haaaa;
            14'h0a03: oData <= 16'h80aa;
            14'h0a04: oData <= 16'ha8aa;
            14'h0a05: oData <= 16'h002a;
            14'h0a06: oData <= 16'hfa80;
            14'h0a07: oData <= 16'hffff;
            14'h0a08: oData <= 16'haffa;
            14'h0a09: oData <= 16'hfffe;
            14'h0a0a: oData <= 16'hffff;
            14'h0a0b: oData <= 16'haaab;
            14'h0a0c: oData <= 16'haaaa;
            14'h0a0d: oData <= 16'hfffa;
            14'h0a0e: oData <= 16'habfa;
            14'h0a0f: oData <= 16'h000a;
            14'h0a10: oData <= 16'h0000;
            14'h0a11: oData <= 16'h0000;
            14'h0a12: oData <= 16'h0000;
            14'h0a13: oData <= 16'h0000;
            14'h0a14: oData <= 16'h0000;
            14'h0a15: oData <= 16'ha000;
            14'h0a16: oData <= 16'h802a;
            14'h0a17: oData <= 16'h00aa;
            14'h0a18: oData <= 16'haaaa;
            14'h0a19: oData <= 16'h002a;
            14'h0a1a: oData <= 16'hfea0;
            14'h0a1b: oData <= 16'hafff;
            14'h0a1c: oData <= 16'hfaff;
            14'h0a1d: oData <= 16'haaff;
            14'h0a1e: oData <= 16'hfaaa;
            14'h0a1f: oData <= 16'hffff;
            14'h0a20: oData <= 16'hffff;
            14'h0a21: oData <= 16'hffff;
            14'h0a22: oData <= 16'hbffb;
            14'h0a23: oData <= 16'h002a;
            14'h0a24: oData <= 16'h0000;
            14'h0a25: oData <= 16'h0000;
            14'h0a26: oData <= 16'h0000;
            14'h0a27: oData <= 16'h0000;
            14'h0a28: oData <= 16'h0000;
            14'h0a29: oData <= 16'ha000;
            14'h0a2a: oData <= 16'h000a;
            14'h0a2b: oData <= 16'h02aa;
            14'h0a2c: oData <= 16'haaaa;
            14'h0a2d: oData <= 16'h000a;
            14'h0a2e: oData <= 16'hffa8;
            14'h0a2f: oData <= 16'hfbff;
            14'h0a30: oData <= 16'hffaf;
            14'h0a31: oData <= 16'hffaa;
            14'h0a32: oData <= 16'hebff;
            14'h0a33: oData <= 16'hffff;
            14'h0a34: oData <= 16'hffff;
            14'h0a35: oData <= 16'hfaab;
            14'h0a36: oData <= 16'hffff;
            14'h0a37: oData <= 16'h00ab;
            14'h0a38: oData <= 16'h0000;
            14'h0a39: oData <= 16'h0000;
            14'h0a3a: oData <= 16'h0000;
            14'h0a3b: oData <= 16'h0000;
            14'h0a3c: oData <= 16'h0000;
            14'h0a3d: oData <= 16'ha800;
            14'h0a3e: oData <= 16'h000a;
            14'h0a3f: oData <= 16'h02aa;
            14'h0a40: oData <= 16'haaa8;
            14'h0a41: oData <= 16'h0000;
            14'h0a42: oData <= 16'hffe8;
            14'h0a43: oData <= 16'hfebf;
            14'h0a44: oData <= 16'habfa;
            14'h0a45: oData <= 16'hffff;
            14'h0a46: oData <= 16'hfebf;
            14'h0a47: oData <= 16'hffff;
            14'h0a48: oData <= 16'haaff;
            14'h0a49: oData <= 16'hebfe;
            14'h0a4a: oData <= 16'hffff;
            14'h0a4b: oData <= 16'h02af;
            14'h0a4c: oData <= 16'h0000;
            14'h0a4d: oData <= 16'h0000;
            14'h0a4e: oData <= 16'h0000;
            14'h0a4f: oData <= 16'h0000;
            14'h0a50: oData <= 16'h0000;
            14'h0a51: oData <= 16'ha800;
            14'h0a52: oData <= 16'h000a;
            14'h0a53: oData <= 16'h02a8;
            14'h0a54: oData <= 16'h2aa0;
            14'h0a55: oData <= 16'h0000;
            14'h0a56: oData <= 16'hffea;
            14'h0a57: oData <= 16'hbfef;
            14'h0a58: oData <= 16'hfebf;
            14'h0a59: oData <= 16'hffff;
            14'h0a5a: oData <= 16'hfaff;
            14'h0a5b: oData <= 16'hffff;
            14'h0a5c: oData <= 16'hffab;
            14'h0a5d: oData <= 16'hbfff;
            14'h0a5e: oData <= 16'hfffe;
            14'h0a5f: oData <= 16'h02bf;
            14'h0a60: oData <= 16'h0000;
            14'h0a61: oData <= 16'h0000;
            14'h0a62: oData <= 16'h0000;
            14'h0a63: oData <= 16'h0000;
            14'h0a64: oData <= 16'h0000;
            14'h0a65: oData <= 16'ha800;
            14'h0a66: oData <= 16'h000a;
            14'h0a67: oData <= 16'h02a8;
            14'h0a68: oData <= 16'h2aa0;
            14'h0a69: oData <= 16'h0000;
            14'h0a6a: oData <= 16'hfffa;
            14'h0a6b: oData <= 16'heffb;
            14'h0a6c: oData <= 16'hffef;
            14'h0a6d: oData <= 16'hffff;
            14'h0a6e: oData <= 16'hfbff;
            14'h0a6f: oData <= 16'hffff;
            14'h0a70: oData <= 16'hfffb;
            14'h0a71: oData <= 16'hffff;
            14'h0a72: oData <= 16'hfffb;
            14'h0a73: oData <= 16'h02bf;
            14'h0a74: oData <= 16'h0000;
            14'h0a75: oData <= 16'h0000;
            14'h0a76: oData <= 16'h0000;
            14'h0a77: oData <= 16'h0000;
            14'h0a78: oData <= 16'h00a8;
            14'h0a79: oData <= 16'ha800;
            14'h0a7a: oData <= 16'h000a;
            14'h0a7b: oData <= 16'h02a8;
            14'h0a7c: oData <= 16'h0a80;
            14'h0a7d: oData <= 16'h0000;
            14'h0a7e: oData <= 16'hfffa;
            14'h0a7f: oData <= 16'hfbff;
            14'h0a80: oData <= 16'hfffb;
            14'h0a81: oData <= 16'hffff;
            14'h0a82: oData <= 16'hebff;
            14'h0a83: oData <= 16'hffff;
            14'h0a84: oData <= 16'hfeff;
            14'h0a85: oData <= 16'hffff;
            14'h0a86: oData <= 16'hfffb;
            14'h0a87: oData <= 16'h02bf;
            14'h0a88: oData <= 16'h0000;
            14'h0a89: oData <= 16'h0000;
            14'h0a8a: oData <= 16'h0000;
            14'h0a8b: oData <= 16'h0000;
            14'h0a8c: oData <= 16'h02aa;
            14'h0a8d: oData <= 16'ha000;
            14'h0a8e: oData <= 16'h000a;
            14'h0a8f: oData <= 16'h02a8;
            14'h0a90: oData <= 16'h0000;
            14'h0a91: oData <= 16'h8000;
            14'h0a92: oData <= 16'hfffa;
            14'h0a93: oData <= 16'hfeff;
            14'h0a94: oData <= 16'hfffe;
            14'h0a95: oData <= 16'hffff;
            14'h0a96: oData <= 16'hefff;
            14'h0a97: oData <= 16'hffff;
            14'h0a98: oData <= 16'hffbf;
            14'h0a99: oData <= 16'hffff;
            14'h0a9a: oData <= 16'hffef;
            14'h0a9b: oData <= 16'h02bf;
            14'h0a9c: oData <= 16'h0000;
            14'h0a9d: oData <= 16'h0000;
            14'h0a9e: oData <= 16'h0000;
            14'h0a9f: oData <= 16'h0000;
            14'h0aa0: oData <= 16'h02aa;
            14'h0aa1: oData <= 16'ha000;
            14'h0aa2: oData <= 16'h002a;
            14'h0aa3: oData <= 16'h02a8;
            14'h0aa4: oData <= 16'h0000;
            14'h0aa5: oData <= 16'h8000;
            14'h0aa6: oData <= 16'hfffe;
            14'h0aa7: oData <= 16'hbfff;
            14'h0aa8: oData <= 16'hffff;
            14'h0aa9: oData <= 16'heaaa;
            14'h0aaa: oData <= 16'hefff;
            14'h0aab: oData <= 16'hffff;
            14'h0aac: oData <= 16'hffef;
            14'h0aad: oData <= 16'hffff;
            14'h0aae: oData <= 16'hffef;
            14'h0aaf: oData <= 16'h0abf;
            14'h0ab0: oData <= 16'h0000;
            14'h0ab1: oData <= 16'h0000;
            14'h0ab2: oData <= 16'h0000;
            14'h0ab3: oData <= 16'h0000;
            14'h0ab4: oData <= 16'h0aaa;
            14'h0ab5: oData <= 16'ha000;
            14'h0ab6: oData <= 16'h00aa;
            14'h0ab7: oData <= 16'h02aa;
            14'h0ab8: oData <= 16'h0000;
            14'h0ab9: oData <= 16'ha000;
            14'h0aba: oData <= 16'hfffe;
            14'h0abb: oData <= 16'hffff;
            14'h0abc: oData <= 16'haaff;
            14'h0abd: oData <= 16'haaaa;
            14'h0abe: oData <= 16'heffa;
            14'h0abf: oData <= 16'hffff;
            14'h0ac0: oData <= 16'hffef;
            14'h0ac1: oData <= 16'hffff;
            14'h0ac2: oData <= 16'hffff;
            14'h0ac3: oData <= 16'h0aff;
            14'h0ac4: oData <= 16'h0000;
            14'h0ac5: oData <= 16'h0000;
            14'h0ac6: oData <= 16'h0000;
            14'h0ac7: oData <= 16'h0000;
            14'h0ac8: oData <= 16'h0aa8;
            14'h0ac9: oData <= 16'h8000;
            14'h0aca: oData <= 16'haaaa;
            14'h0acb: oData <= 16'h02aa;
            14'h0acc: oData <= 16'h0000;
            14'h0acd: oData <= 16'ha800;
            14'h0ace: oData <= 16'hffff;
            14'h0acf: oData <= 16'hffff;
            14'h0ad0: oData <= 16'haaaf;
            14'h0ad1: oData <= 16'haeaa;
            14'h0ad2: oData <= 16'hffaa;
            14'h0ad3: oData <= 16'hffff;
            14'h0ad4: oData <= 16'hffef;
            14'h0ad5: oData <= 16'hffff;
            14'h0ad6: oData <= 16'hffff;
            14'h0ad7: oData <= 16'h0aff;
            14'h0ad8: oData <= 16'h0000;
            14'h0ad9: oData <= 16'h0000;
            14'h0ada: oData <= 16'h0000;
            14'h0adb: oData <= 16'h0000;
            14'h0adc: oData <= 16'h2aa8;
            14'h0add: oData <= 16'h0000;
            14'h0ade: oData <= 16'haaaa;
            14'h0adf: oData <= 16'h00aa;
            14'h0ae0: oData <= 16'h0000;
            14'h0ae1: oData <= 16'hea00;
            14'h0ae2: oData <= 16'hffff;
            14'h0ae3: oData <= 16'hffff;
            14'h0ae4: oData <= 16'haaab;
            14'h0ae5: oData <= 16'hfeaa;
            14'h0ae6: oData <= 16'hfeab;
            14'h0ae7: oData <= 16'hffff;
            14'h0ae8: oData <= 16'hafef;
            14'h0ae9: oData <= 16'haaaa;
            14'h0aea: oData <= 16'hffff;
            14'h0aeb: oData <= 16'h2aff;
            14'h0aec: oData <= 16'h0000;
            14'h0aed: oData <= 16'h0000;
            14'h0aee: oData <= 16'h0000;
            14'h0aef: oData <= 16'h0000;
            14'h0af0: oData <= 16'h2aa0;
            14'h0af1: oData <= 16'h0000;
            14'h0af2: oData <= 16'haaaa;
            14'h0af3: oData <= 16'h00aa;
            14'h0af4: oData <= 16'h0000;
            14'h0af5: oData <= 16'haa80;
            14'h0af6: oData <= 16'hffaa;
            14'h0af7: oData <= 16'hfaff;
            14'h0af8: oData <= 16'habea;
            14'h0af9: oData <= 16'hfeaa;
            14'h0afa: oData <= 16'heabf;
            14'h0afb: oData <= 16'hffff;
            14'h0afc: oData <= 16'haaff;
            14'h0afd: oData <= 16'hbffa;
            14'h0afe: oData <= 16'hfffa;
            14'h0aff: oData <= 16'habff;
            14'h0b00: oData <= 16'h0002;
            14'h0b01: oData <= 16'h0000;
            14'h0b02: oData <= 16'h0000;
            14'h0b03: oData <= 16'h0000;
            14'h0b04: oData <= 16'h2aa0;
            14'h0b05: oData <= 16'h0000;
            14'h0b06: oData <= 16'haaa8;
            14'h0b07: oData <= 16'h002a;
            14'h0b08: oData <= 16'h0000;
            14'h0b09: oData <= 16'hfaa0;
            14'h0b0a: oData <= 16'hffff;
            14'h0b0b: oData <= 16'hbfaf;
            14'h0b0c: oData <= 16'haaaa;
            14'h0b0d: oData <= 16'heaaa;
            14'h0b0e: oData <= 16'heaff;
            14'h0b0f: oData <= 16'hffff;
            14'h0b10: oData <= 16'haabf;
            14'h0b11: oData <= 16'haaaa;
            14'h0b12: oData <= 16'hfefa;
            14'h0b13: oData <= 16'hafff;
            14'h0b14: oData <= 16'h000a;
            14'h0b15: oData <= 16'h0000;
            14'h0b16: oData <= 16'h0000;
            14'h0b17: oData <= 16'h0000;
            14'h0b18: oData <= 16'haaa0;
            14'h0b19: oData <= 16'h0000;
            14'h0b1a: oData <= 16'h0000;
            14'h0b1b: oData <= 16'h0000;
            14'h0b1c: oData <= 16'h0000;
            14'h0b1d: oData <= 16'haba8;
            14'h0b1e: oData <= 16'hfaaa;
            14'h0b1f: oData <= 16'hbebf;
            14'h0b20: oData <= 16'haaaa;
            14'h0b21: oData <= 16'haaaa;
            14'h0b22: oData <= 16'habfe;
            14'h0b23: oData <= 16'hbfff;
            14'h0b24: oData <= 16'haaae;
            14'h0b25: oData <= 16'haaaa;
            14'h0b26: oData <= 16'hbaba;
            14'h0b27: oData <= 16'hfeaa;
            14'h0b28: oData <= 16'h002a;
            14'h0b29: oData <= 16'h0000;
            14'h0b2a: oData <= 16'h0000;
            14'h0b2b: oData <= 16'h0000;
            14'h0b2c: oData <= 16'haa80;
            14'h0b2d: oData <= 16'h0000;
            14'h0b2e: oData <= 16'h0000;
            14'h0b2f: oData <= 16'h0000;
            14'h0b30: oData <= 16'h0000;
            14'h0b31: oData <= 16'hfeea;
            14'h0b32: oData <= 16'hffff;
            14'h0b33: oData <= 16'hebff;
            14'h0b34: oData <= 16'hffeb;
            14'h0b35: oData <= 16'hafff;
            14'h0b36: oData <= 16'heaaa;
            14'h0b37: oData <= 16'hafff;
            14'h0b38: oData <= 16'haaaa;
            14'h0b39: oData <= 16'hffea;
            14'h0b3a: oData <= 16'hefff;
            14'h0b3b: oData <= 16'hfbff;
            14'h0b3c: oData <= 16'h002b;
            14'h0b3d: oData <= 16'h0000;
            14'h0b3e: oData <= 16'h0000;
            14'h0b3f: oData <= 16'h0000;
            14'h0b40: oData <= 16'haa80;
            14'h0b41: oData <= 16'ha000;
            14'h0b42: oData <= 16'h0002;
            14'h0b43: oData <= 16'h0000;
            14'h0b44: oData <= 16'h8000;
            14'h0b45: oData <= 16'hffba;
            14'h0b46: oData <= 16'haaab;
            14'h0b47: oData <= 16'hfbfe;
            14'h0b48: oData <= 16'hffff;
            14'h0b49: oData <= 16'hffea;
            14'h0b4a: oData <= 16'heaaa;
            14'h0b4b: oData <= 16'hffff;
            14'h0b4c: oData <= 16'hfaaa;
            14'h0b4d: oData <= 16'hffff;
            14'h0b4e: oData <= 16'hffff;
            14'h0b4f: oData <= 16'hefaf;
            14'h0b50: oData <= 16'h00ab;
            14'h0b51: oData <= 16'h0000;
            14'h0b52: oData <= 16'h0000;
            14'h0b53: oData <= 16'h0000;
            14'h0b54: oData <= 16'haa80;
            14'h0b55: oData <= 16'ha802;
            14'h0b56: oData <= 16'h000a;
            14'h0b57: oData <= 16'h0000;
            14'h0b58: oData <= 16'ha000;
            14'h0b59: oData <= 16'hbfee;
            14'h0b5a: oData <= 16'haaaa;
            14'h0b5b: oData <= 16'hffaa;
            14'h0b5c: oData <= 16'hbfff;
            14'h0b5d: oData <= 16'hfffa;
            14'h0b5e: oData <= 16'hfebf;
            14'h0b5f: oData <= 16'hffff;
            14'h0b60: oData <= 16'hffaf;
            14'h0b61: oData <= 16'hffff;
            14'h0b62: oData <= 16'hffff;
            14'h0b63: oData <= 16'hbeff;
            14'h0b64: oData <= 16'h00ae;
            14'h0b65: oData <= 16'h0000;
            14'h0b66: oData <= 16'h0000;
            14'h0b67: oData <= 16'h0000;
            14'h0b68: oData <= 16'haa00;
            14'h0b69: oData <= 16'haa82;
            14'h0b6a: oData <= 16'h000a;
            14'h0b6b: oData <= 16'h0000;
            14'h0b6c: oData <= 16'ha000;
            14'h0b6d: oData <= 16'haffb;
            14'h0b6e: oData <= 16'hfffa;
            14'h0b6f: oData <= 16'hfaaa;
            14'h0b70: oData <= 16'habff;
            14'h0b71: oData <= 16'hfffe;
            14'h0b72: oData <= 16'hffff;
            14'h0b73: oData <= 16'hffff;
            14'h0b74: oData <= 16'hffaf;
            14'h0b75: oData <= 16'hffff;
            14'h0b76: oData <= 16'haaff;
            14'h0b77: oData <= 16'hfbfa;
            14'h0b78: oData <= 16'h00ae;
            14'h0b79: oData <= 16'h0000;
            14'h0b7a: oData <= 16'h0000;
            14'h0b7b: oData <= 16'h0000;
            14'h0b7c: oData <= 16'haa00;
            14'h0b7d: oData <= 16'haaaa;
            14'h0b7e: oData <= 16'h000a;
            14'h0b7f: oData <= 16'h0000;
            14'h0b80: oData <= 16'ha800;
            14'h0b81: oData <= 16'haffb;
            14'h0b82: oData <= 16'hefff;
            14'h0b83: oData <= 16'haaaf;
            14'h0b84: oData <= 16'haaaa;
            14'h0b85: oData <= 16'hffff;
            14'h0b86: oData <= 16'hffff;
            14'h0b87: oData <= 16'hffff;
            14'h0b88: oData <= 16'hffaf;
            14'h0b89: oData <= 16'hffff;
            14'h0b8a: oData <= 16'haabf;
            14'h0b8b: oData <= 16'hfbaa;
            14'h0b8c: oData <= 16'h00ab;
            14'h0b8d: oData <= 16'h0000;
            14'h0b8e: oData <= 16'h0000;
            14'h0b8f: oData <= 16'h0000;
            14'h0b90: oData <= 16'haa00;
            14'h0b91: oData <= 16'haaaa;
            14'h0b92: oData <= 16'h0002;
            14'h0b93: oData <= 16'h0000;
            14'h0b94: oData <= 16'he800;
            14'h0b95: oData <= 16'habfb;
            14'h0b96: oData <= 16'hebff;
            14'h0b97: oData <= 16'habff;
            14'h0b98: oData <= 16'hfaaa;
            14'h0b99: oData <= 16'hffff;
            14'h0b9a: oData <= 16'hffff;
            14'h0b9b: oData <= 16'hffff;
            14'h0b9c: oData <= 16'hffaf;
            14'h0b9d: oData <= 16'hfaff;
            14'h0b9e: oData <= 16'hfeab;
            14'h0b9f: oData <= 16'hfbab;
            14'h0ba0: oData <= 16'h00ab;
            14'h0ba1: oData <= 16'h0000;
            14'h0ba2: oData <= 16'h0000;
            14'h0ba3: oData <= 16'h0000;
            14'h0ba4: oData <= 16'ha800;
            14'h0ba5: oData <= 16'haaaa;
            14'h0ba6: oData <= 16'h0000;
            14'h0ba7: oData <= 16'h0000;
            14'h0ba8: oData <= 16'hea00;
            14'h0ba9: oData <= 16'hebfb;
            14'h0baa: oData <= 16'hebff;
            14'h0bab: oData <= 16'hffff;
            14'h0bac: oData <= 16'hffff;
            14'h0bad: oData <= 16'hffff;
            14'h0bae: oData <= 16'hffff;
            14'h0baf: oData <= 16'hffff;
            14'h0bb0: oData <= 16'hffaf;
            14'h0bb1: oData <= 16'haaff;
            14'h0bb2: oData <= 16'hffaa;
            14'h0bb3: oData <= 16'hfbbf;
            14'h0bb4: oData <= 16'h00ab;
            14'h0bb5: oData <= 16'h0000;
            14'h0bb6: oData <= 16'h0000;
            14'h0bb7: oData <= 16'h0000;
            14'h0bb8: oData <= 16'ha800;
            14'h0bb9: oData <= 16'h0aaa;
            14'h0bba: oData <= 16'h0000;
            14'h0bbb: oData <= 16'h0000;
            14'h0bbc: oData <= 16'hfa00;
            14'h0bbd: oData <= 16'heafb;
            14'h0bbe: oData <= 16'habff;
            14'h0bbf: oData <= 16'hfffe;
            14'h0bc0: oData <= 16'hffff;
            14'h0bc1: oData <= 16'hffff;
            14'h0bc2: oData <= 16'hffff;
            14'h0bc3: oData <= 16'hffff;
            14'h0bc4: oData <= 16'hfaaf;
            14'h0bc5: oData <= 16'habff;
            14'h0bc6: oData <= 16'hefea;
            14'h0bc7: oData <= 16'hefff;
            14'h0bc8: oData <= 16'h00ab;
            14'h0bc9: oData <= 16'h0000;
            14'h0bca: oData <= 16'h0000;
            14'h0bcb: oData <= 16'h0000;
            14'h0bcc: oData <= 16'ha800;
            14'h0bcd: oData <= 16'h00aa;
            14'h0bce: oData <= 16'h0000;
            14'h0bcf: oData <= 16'h0000;
            14'h0bd0: oData <= 16'hfa00;
            14'h0bd1: oData <= 16'hfafb;
            14'h0bd2: oData <= 16'haaff;
            14'h0bd3: oData <= 16'hffea;
            14'h0bd4: oData <= 16'hffff;
            14'h0bd5: oData <= 16'hbfff;
            14'h0bd6: oData <= 16'hfaaf;
            14'h0bd7: oData <= 16'hffff;
            14'h0bd8: oData <= 16'heabf;
            14'h0bd9: oData <= 16'hffff;
            14'h0bda: oData <= 16'hebff;
            14'h0bdb: oData <= 16'hefff;
            14'h0bdc: oData <= 16'h00ab;
            14'h0bdd: oData <= 16'h0000;
            14'h0bde: oData <= 16'h0000;
            14'h0bdf: oData <= 16'h0000;
            14'h0be0: oData <= 16'ha000;
            14'h0be1: oData <= 16'h000a;
            14'h0be2: oData <= 16'h0000;
            14'h0be3: oData <= 16'h0000;
            14'h0be4: oData <= 16'hfa00;
            14'h0be5: oData <= 16'hfafb;
            14'h0be6: oData <= 16'hfaaf;
            14'h0be7: oData <= 16'hfeaa;
            14'h0be8: oData <= 16'hffff;
            14'h0be9: oData <= 16'hbfff;
            14'h0bea: oData <= 16'heaab;
            14'h0beb: oData <= 16'hffff;
            14'h0bec: oData <= 16'habff;
            14'h0bed: oData <= 16'hfffe;
            14'h0bee: oData <= 16'hebff;
            14'h0bef: oData <= 16'hefff;
            14'h0bf0: oData <= 16'h00ab;
            14'h0bf1: oData <= 16'h0000;
            14'h0bf2: oData <= 16'h0000;
            14'h0bf3: oData <= 16'h0000;
            14'h0bf4: oData <= 16'h0000;
            14'h0bf5: oData <= 16'h0000;
            14'h0bf6: oData <= 16'h0000;
            14'h0bf7: oData <= 16'h0000;
            14'h0bf8: oData <= 16'hea00;
            14'h0bf9: oData <= 16'hfafb;
            14'h0bfa: oData <= 16'hfaaa;
            14'h0bfb: oData <= 16'heaaf;
            14'h0bfc: oData <= 16'hbfff;
            14'h0bfd: oData <= 16'heaaa;
            14'h0bfe: oData <= 16'hffea;
            14'h0bff: oData <= 16'hffff;
            14'h0c00: oData <= 16'hafff;
            14'h0c01: oData <= 16'hfffa;
            14'h0c02: oData <= 16'hebff;
            14'h0c03: oData <= 16'hfbff;
            14'h0c04: oData <= 16'h00ae;
            14'h0c05: oData <= 16'h0000;
            14'h0c06: oData <= 16'h0000;
            14'h0c07: oData <= 16'h0000;
            14'h0c08: oData <= 16'h0000;
            14'h0c09: oData <= 16'h0000;
            14'h0c0a: oData <= 16'h0000;
            14'h0c0b: oData <= 16'h0000;
            14'h0c0c: oData <= 16'he800;
            14'h0c0d: oData <= 16'heafb;
            14'h0c0e: oData <= 16'heaea;
            14'h0c0f: oData <= 16'haaff;
            14'h0c10: oData <= 16'hbffa;
            14'h0c11: oData <= 16'hffff;
            14'h0c12: oData <= 16'hfffa;
            14'h0c13: oData <= 16'hffff;
            14'h0c14: oData <= 16'hafff;
            14'h0c15: oData <= 16'hffea;
            14'h0c16: oData <= 16'habff;
            14'h0c17: oData <= 16'hfebe;
            14'h0c18: oData <= 16'h00aa;
            14'h0c19: oData <= 16'h0000;
            14'h0c1a: oData <= 16'h0000;
            14'h0c1b: oData <= 16'h0000;
            14'h0c1c: oData <= 16'h0000;
            14'h0c1d: oData <= 16'h0000;
            14'h0c1e: oData <= 16'h0000;
            14'h0c1f: oData <= 16'h0000;
            14'h0c20: oData <= 16'he800;
            14'h0c21: oData <= 16'hebfb;
            14'h0c22: oData <= 16'hebff;
            14'h0c23: oData <= 16'hafff;
            14'h0c24: oData <= 16'hffaa;
            14'h0c25: oData <= 16'hffff;
            14'h0c26: oData <= 16'habfa;
            14'h0c27: oData <= 16'hffaa;
            14'h0c28: oData <= 16'habff;
            14'h0c29: oData <= 16'hfeba;
            14'h0c2a: oData <= 16'habff;
            14'h0c2b: oData <= 16'hbffe;
            14'h0c2c: oData <= 16'h002b;
            14'h0c2d: oData <= 16'h0000;
            14'h0c2e: oData <= 16'h0000;
            14'h0c2f: oData <= 16'h0000;
            14'h0c30: oData <= 16'h0000;
            14'h0c31: oData <= 16'h0000;
            14'h0c32: oData <= 16'h0000;
            14'h0c33: oData <= 16'h0000;
            14'h0c34: oData <= 16'he800;
            14'h0c35: oData <= 16'habef;
            14'h0c36: oData <= 16'habff;
            14'h0c37: oData <= 16'hffff;
            14'h0c38: oData <= 16'heaaa;
            14'h0c39: oData <= 16'hffff;
            14'h0c3a: oData <= 16'habea;
            14'h0c3b: oData <= 16'hffaa;
            14'h0c3c: oData <= 16'hebff;
            14'h0c3d: oData <= 16'hebfa;
            14'h0c3e: oData <= 16'haaff;
            14'h0c3f: oData <= 16'heafe;
            14'h0c40: oData <= 16'h002b;
            14'h0c41: oData <= 16'h0000;
            14'h0c42: oData <= 16'h0000;
            14'h0c43: oData <= 16'h0000;
            14'h0c44: oData <= 16'h0000;
            14'h0c45: oData <= 16'h0000;
            14'h0c46: oData <= 16'h0000;
            14'h0c47: oData <= 16'h0000;
            14'h0c48: oData <= 16'ha800;
            14'h0c49: oData <= 16'hafef;
            14'h0c4a: oData <= 16'habff;
            14'h0c4b: oData <= 16'hfffe;
            14'h0c4c: oData <= 16'haaba;
            14'h0c4d: oData <= 16'hffea;
            14'h0c4e: oData <= 16'hfbab;
            14'h0c4f: oData <= 16'hffff;
            14'h0c50: oData <= 16'heaff;
            14'h0c51: oData <= 16'hbfff;
            14'h0c52: oData <= 16'hbabf;
            14'h0c53: oData <= 16'hffbe;
            14'h0c54: oData <= 16'h002a;
            14'h0c55: oData <= 16'h0000;
            14'h0c56: oData <= 16'h0000;
            14'h0c57: oData <= 16'h0000;
            14'h0c58: oData <= 16'h0000;
            14'h0c59: oData <= 16'h0000;
            14'h0c5a: oData <= 16'h0000;
            14'h0c5b: oData <= 16'h0000;
            14'h0c5c: oData <= 16'ha000;
            14'h0c5d: oData <= 16'hffbe;
            14'h0c5e: oData <= 16'habff;
            14'h0c5f: oData <= 16'hffea;
            14'h0c60: oData <= 16'haffa;
            14'h0c61: oData <= 16'hfaaa;
            14'h0c62: oData <= 16'hffef;
            14'h0c63: oData <= 16'hbfff;
            14'h0c64: oData <= 16'hfaae;
            14'h0c65: oData <= 16'hffff;
            14'h0c66: oData <= 16'haaaf;
            14'h0c67: oData <= 16'hbffe;
            14'h0c68: oData <= 16'h000a;
            14'h0c69: oData <= 16'h0000;
            14'h0c6a: oData <= 16'h0000;
            14'h0c6b: oData <= 16'h0000;
            14'h0c6c: oData <= 16'h0000;
            14'h0c6d: oData <= 16'h0000;
            14'h0c6e: oData <= 16'h0000;
            14'h0c6f: oData <= 16'h0000;
            14'h0c70: oData <= 16'h8000;
            14'h0c71: oData <= 16'hfafe;
            14'h0c72: oData <= 16'hafff;
            14'h0c73: oData <= 16'hfeaa;
            14'h0c74: oData <= 16'hfffa;
            14'h0c75: oData <= 16'haaaf;
            14'h0c76: oData <= 16'hfffe;
            14'h0c77: oData <= 16'hbfff;
            14'h0c78: oData <= 16'hfeaa;
            14'h0c79: oData <= 16'hffff;
            14'h0c7a: oData <= 16'habaa;
            14'h0c7b: oData <= 16'hbffa;
            14'h0c7c: oData <= 16'h0002;
            14'h0c7d: oData <= 16'h0000;
            14'h0c7e: oData <= 16'h0000;
            14'h0c7f: oData <= 16'h0000;
            14'h0c80: oData <= 16'h0000;
            14'h0c81: oData <= 16'h0000;
            14'h0c82: oData <= 16'h0000;
            14'h0c83: oData <= 16'h0000;
            14'h0c84: oData <= 16'h8000;
            14'h0c85: oData <= 16'haffa;
            14'h0c86: oData <= 16'hbfff;
            14'h0c87: oData <= 16'heaaa;
            14'h0c88: oData <= 16'hffea;
            14'h0c89: oData <= 16'habff;
            14'h0c8a: oData <= 16'hfeaa;
            14'h0c8b: oData <= 16'hffff;
            14'h0c8c: oData <= 16'hffea;
            14'h0c8d: oData <= 16'hafff;
            14'h0c8e: oData <= 16'hebaa;
            14'h0c8f: oData <= 16'haffa;
            14'h0c90: oData <= 16'h0002;
            14'h0c91: oData <= 16'h0000;
            14'h0c92: oData <= 16'h0000;
            14'h0c93: oData <= 16'h0000;
            14'h0c94: oData <= 16'h0000;
            14'h0c95: oData <= 16'h0000;
            14'h0c96: oData <= 16'h0000;
            14'h0c97: oData <= 16'h0000;
            14'h0c98: oData <= 16'h0000;
            14'h0c99: oData <= 16'hfeaa;
            14'h0c9a: oData <= 16'hffff;
            14'h0c9b: oData <= 16'haaba;
            14'h0c9c: oData <= 16'hffaa;
            14'h0c9d: oData <= 16'hafff;
            14'h0c9e: oData <= 16'haaaa;
            14'h0c9f: oData <= 16'hffea;
            14'h0ca0: oData <= 16'hffff;
            14'h0ca1: oData <= 16'haabf;
            14'h0ca2: oData <= 16'habae;
            14'h0ca3: oData <= 16'haffa;
            14'h0ca4: oData <= 16'h0000;
            14'h0ca5: oData <= 16'h0000;
            14'h0ca6: oData <= 16'h0000;
            14'h0ca7: oData <= 16'h0000;
            14'h0ca8: oData <= 16'h0000;
            14'h0ca9: oData <= 16'h0000;
            14'h0caa: oData <= 16'h0000;
            14'h0cab: oData <= 16'h0000;
            14'h0cac: oData <= 16'h0000;
            14'h0cad: oData <= 16'hfba8;
            14'h0cae: oData <= 16'hffff;
            14'h0caf: oData <= 16'hafea;
            14'h0cb0: oData <= 16'hfeaa;
            14'h0cb1: oData <= 16'hafff;
            14'h0cb2: oData <= 16'haaff;
            14'h0cb3: oData <= 16'haaaa;
            14'h0cb4: oData <= 16'haaaa;
            14'h0cb5: oData <= 16'heaaa;
            14'h0cb6: oData <= 16'hafaf;
            14'h0cb7: oData <= 16'haffa;
            14'h0cb8: oData <= 16'h0000;
            14'h0cb9: oData <= 16'h0000;
            14'h0cba: oData <= 16'h0000;
            14'h0cbb: oData <= 16'h0000;
            14'h0cbc: oData <= 16'h0000;
            14'h0cbd: oData <= 16'h0000;
            14'h0cbe: oData <= 16'h0000;
            14'h0cbf: oData <= 16'h0000;
            14'h0cc0: oData <= 16'h0000;
            14'h0cc1: oData <= 16'hfea0;
            14'h0cc2: oData <= 16'hffff;
            14'h0cc3: oData <= 16'hffab;
            14'h0cc4: oData <= 16'haaaa;
            14'h0cc5: oData <= 16'hafff;
            14'h0cc6: oData <= 16'hffff;
            14'h0cc7: oData <= 16'haaaf;
            14'h0cc8: oData <= 16'haaaa;
            14'h0cc9: oData <= 16'hfaaa;
            14'h0cca: oData <= 16'hafaf;
            14'h0ccb: oData <= 16'haffa;
            14'h0ccc: oData <= 16'h0000;
            14'h0ccd: oData <= 16'h0000;
            14'h0cce: oData <= 16'h0000;
            14'h0ccf: oData <= 16'h0000;
            14'h0cd0: oData <= 16'h0000;
            14'h0cd1: oData <= 16'h0000;
            14'h0cd2: oData <= 16'h0000;
            14'h0cd3: oData <= 16'h0000;
            14'h0cd4: oData <= 16'h0000;
            14'h0cd5: oData <= 16'hfa80;
            14'h0cd6: oData <= 16'hffff;
            14'h0cd7: oData <= 16'hffaf;
            14'h0cd8: oData <= 16'haaaa;
            14'h0cd9: oData <= 16'habea;
            14'h0cda: oData <= 16'hffff;
            14'h0cdb: oData <= 16'hffaf;
            14'h0cdc: oData <= 16'hfebf;
            14'h0cdd: oData <= 16'heaff;
            14'h0cde: oData <= 16'hafaf;
            14'h0cdf: oData <= 16'haffa;
            14'h0ce0: oData <= 16'h0000;
            14'h0ce1: oData <= 16'h0000;
            14'h0ce2: oData <= 16'h0000;
            14'h0ce3: oData <= 16'h0000;
            14'h0ce4: oData <= 16'h0000;
            14'h0ce5: oData <= 16'h0000;
            14'h0ce6: oData <= 16'h0000;
            14'h0ce7: oData <= 16'h0000;
            14'h0ce8: oData <= 16'h0000;
            14'h0ce9: oData <= 16'hea00;
            14'h0cea: oData <= 16'hffff;
            14'h0ceb: oData <= 16'hfeaf;
            14'h0cec: oData <= 16'haafa;
            14'h0ced: oData <= 16'heaaa;
            14'h0cee: oData <= 16'hffff;
            14'h0cef: oData <= 16'hffaf;
            14'h0cf0: oData <= 16'hfebf;
            14'h0cf1: oData <= 16'hebff;
            14'h0cf2: oData <= 16'habaf;
            14'h0cf3: oData <= 16'haffa;
            14'h0cf4: oData <= 16'h0000;
            14'h0cf5: oData <= 16'h0000;
            14'h0cf6: oData <= 16'h0000;
            14'h0cf7: oData <= 16'h0000;
            14'h0cf8: oData <= 16'h0000;
            14'h0cf9: oData <= 16'h0000;
            14'h0cfa: oData <= 16'h0000;
            14'h0cfb: oData <= 16'h0000;
            14'h0cfc: oData <= 16'h0000;
            14'h0cfd: oData <= 16'ha800;
            14'h0cfe: oData <= 16'hffff;
            14'h0cff: oData <= 16'hfabf;
            14'h0d00: oData <= 16'haffa;
            14'h0d01: oData <= 16'haaaa;
            14'h0d02: oData <= 16'hfffe;
            14'h0d03: oData <= 16'hffaf;
            14'h0d04: oData <= 16'hfebf;
            14'h0d05: oData <= 16'hebff;
            14'h0d06: oData <= 16'haaaf;
            14'h0d07: oData <= 16'haffa;
            14'h0d08: oData <= 16'h0000;
            14'h0d09: oData <= 16'h0000;
            14'h0d0a: oData <= 16'h0000;
            14'h0d0b: oData <= 16'h0000;
            14'h0d0c: oData <= 16'h0000;
            14'h0d0d: oData <= 16'h0000;
            14'h0d0e: oData <= 16'h0000;
            14'h0d0f: oData <= 16'h0000;
            14'h0d10: oData <= 16'h0000;
            14'h0d11: oData <= 16'ha000;
            14'h0d12: oData <= 16'hffff;
            14'h0d13: oData <= 16'heaff;
            14'h0d14: oData <= 16'hfffa;
            14'h0d15: oData <= 16'haaaa;
            14'h0d16: oData <= 16'hfeaa;
            14'h0d17: oData <= 16'hffaf;
            14'h0d18: oData <= 16'hfebf;
            14'h0d19: oData <= 16'haaaf;
            14'h0d1a: oData <= 16'haaaa;
            14'h0d1b: oData <= 16'haffa;
            14'h0d1c: oData <= 16'h0000;
            14'h0d1d: oData <= 16'h0000;
            14'h0d1e: oData <= 16'h0000;
            14'h0d1f: oData <= 16'h0000;
            14'h0d20: oData <= 16'h0000;
            14'h0d21: oData <= 16'h0000;
            14'h0d22: oData <= 16'h0000;
            14'h0d23: oData <= 16'h0000;
            14'h0d24: oData <= 16'h0000;
            14'h0d25: oData <= 16'ha000;
            14'h0d26: oData <= 16'hffff;
            14'h0d27: oData <= 16'habff;
            14'h0d28: oData <= 16'hfffa;
            14'h0d29: oData <= 16'haaff;
            14'h0d2a: oData <= 16'haaaa;
            14'h0d2b: oData <= 16'haaaa;
            14'h0d2c: oData <= 16'haaaa;
            14'h0d2d: oData <= 16'haaaa;
            14'h0d2e: oData <= 16'haaaa;
            14'h0d2f: oData <= 16'haffa;
            14'h0d30: oData <= 16'h0000;
            14'h0d31: oData <= 16'h0000;
            14'h0d32: oData <= 16'h0000;
            14'h0d33: oData <= 16'h0000;
            14'h0d34: oData <= 16'h0000;
            14'h0d35: oData <= 16'h0000;
            14'h0d36: oData <= 16'h0000;
            14'h0d37: oData <= 16'h0000;
            14'h0d38: oData <= 16'h0000;
            14'h0d39: oData <= 16'ha000;
            14'h0d3a: oData <= 16'hfffe;
            14'h0d3b: oData <= 16'hafff;
            14'h0d3c: oData <= 16'hfffe;
            14'h0d3d: oData <= 16'hbaff;
            14'h0d3e: oData <= 16'haaaa;
            14'h0d3f: oData <= 16'haaaa;
            14'h0d40: oData <= 16'haaaa;
            14'h0d41: oData <= 16'haaaa;
            14'h0d42: oData <= 16'haaaa;
            14'h0d43: oData <= 16'haffa;
            14'h0d44: oData <= 16'h0000;
            14'h0d45: oData <= 16'h0000;
            14'h0d46: oData <= 16'h0000;
            14'h0d47: oData <= 16'h0000;
            14'h0d48: oData <= 16'h0000;
            14'h0d49: oData <= 16'h0000;
            14'h0d4a: oData <= 16'h0000;
            14'h0d4b: oData <= 16'h0000;
            14'h0d4c: oData <= 16'h0000;
            14'h0d4d: oData <= 16'h8000;
            14'h0d4e: oData <= 16'hfffe;
            14'h0d4f: oData <= 16'hbfff;
            14'h0d50: oData <= 16'hfffa;
            14'h0d51: oData <= 16'hfaff;
            14'h0d52: oData <= 16'haaaf;
            14'h0d53: oData <= 16'haaaa;
            14'h0d54: oData <= 16'haaaa;
            14'h0d55: oData <= 16'haaaa;
            14'h0d56: oData <= 16'haaaa;
            14'h0d57: oData <= 16'haffa;
            14'h0d58: oData <= 16'h0000;
            14'h0d59: oData <= 16'h0000;
            14'h0d5a: oData <= 16'h0000;
            14'h0d5b: oData <= 16'h0000;
            14'h0d5c: oData <= 16'h0000;
            14'h0d5d: oData <= 16'h0000;
            14'h0d5e: oData <= 16'h0000;
            14'h0d5f: oData <= 16'h0000;
            14'h0d60: oData <= 16'h0000;
            14'h0d61: oData <= 16'h8000;
            14'h0d62: oData <= 16'hfffa;
            14'h0d63: oData <= 16'hffff;
            14'h0d64: oData <= 16'hffea;
            14'h0d65: oData <= 16'hfaff;
            14'h0d66: oData <= 16'habff;
            14'h0d67: oData <= 16'haaaa;
            14'h0d68: oData <= 16'haaaa;
            14'h0d69: oData <= 16'haaaa;
            14'h0d6a: oData <= 16'haaaa;
            14'h0d6b: oData <= 16'haffe;
            14'h0d6c: oData <= 16'h0000;
            14'h0d6d: oData <= 16'h0000;
            14'h0d6e: oData <= 16'h0000;
            14'h0d6f: oData <= 16'h0000;
            14'h0d70: oData <= 16'h0000;
            14'h0d71: oData <= 16'h0000;
            14'h0d72: oData <= 16'h0000;
            14'h0d73: oData <= 16'h0000;
            14'h0d74: oData <= 16'h0000;
            14'h0d75: oData <= 16'h0000;
            14'h0d76: oData <= 16'hffea;
            14'h0d77: oData <= 16'hffff;
            14'h0d78: oData <= 16'hfeab;
            14'h0d79: oData <= 16'hfabf;
            14'h0d7a: oData <= 16'hffff;
            14'h0d7b: oData <= 16'haaaa;
            14'h0d7c: oData <= 16'haaaa;
            14'h0d7d: oData <= 16'haaaa;
            14'h0d7e: oData <= 16'hbaaa;
            14'h0d7f: oData <= 16'haffe;
            14'h0d80: oData <= 16'h0000;
            14'h0d81: oData <= 16'h0000;
            14'h0d82: oData <= 16'h0000;
            14'h0d83: oData <= 16'h0000;
            14'h0d84: oData <= 16'h0000;
            14'h0d85: oData <= 16'h0000;
            14'h0d86: oData <= 16'h0000;
            14'h0d87: oData <= 16'h0000;
            14'h0d88: oData <= 16'h0000;
            14'h0d89: oData <= 16'h02a0;
            14'h0d8a: oData <= 16'hffa8;
            14'h0d8b: oData <= 16'hffff;
            14'h0d8c: oData <= 16'hfaaf;
            14'h0d8d: oData <= 16'hfebf;
            14'h0d8e: oData <= 16'hffff;
            14'h0d8f: oData <= 16'habfa;
            14'h0d90: oData <= 16'haaaa;
            14'h0d91: oData <= 16'haaaa;
            14'h0d92: oData <= 16'hbafa;
            14'h0d93: oData <= 16'haffe;
            14'h0d94: oData <= 16'h0000;
            14'h0d95: oData <= 16'h0000;
            14'h0d96: oData <= 16'h0000;
            14'h0d97: oData <= 16'h0000;
            14'h0d98: oData <= 16'h0000;
            14'h0d99: oData <= 16'h0000;
            14'h0d9a: oData <= 16'h0000;
            14'h0d9b: oData <= 16'h0000;
            14'h0d9c: oData <= 16'h0000;
            14'h0d9d: oData <= 16'h0aa8;
            14'h0d9e: oData <= 16'hfea0;
            14'h0d9f: oData <= 16'hffff;
            14'h0da0: oData <= 16'haaff;
            14'h0da1: oData <= 16'hfebf;
            14'h0da2: oData <= 16'hffff;
            14'h0da3: oData <= 16'hfffa;
            14'h0da4: oData <= 16'hfeaf;
            14'h0da5: oData <= 16'hbfaf;
            14'h0da6: oData <= 16'haebe;
            14'h0da7: oData <= 16'hafff;
            14'h0da8: oData <= 16'h0000;
            14'h0da9: oData <= 16'h0000;
            14'h0daa: oData <= 16'h0000;
            14'h0dab: oData <= 16'h0000;
            14'h0dac: oData <= 16'h0000;
            14'h0dad: oData <= 16'h0000;
            14'h0dae: oData <= 16'h0000;
            14'h0daf: oData <= 16'h0000;
            14'h0db0: oData <= 16'h0000;
            14'h0db1: oData <= 16'h0aa8;
            14'h0db2: oData <= 16'hfaa0;
            14'h0db3: oData <= 16'hffff;
            14'h0db4: oData <= 16'habff;
            14'h0db5: oData <= 16'hfeaa;
            14'h0db6: oData <= 16'hffff;
            14'h0db7: oData <= 16'hfffa;
            14'h0db8: oData <= 16'hffaf;
            14'h0db9: oData <= 16'hafab;
            14'h0dba: oData <= 16'haaae;
            14'h0dbb: oData <= 16'hafff;
            14'h0dbc: oData <= 16'h0000;
            14'h0dbd: oData <= 16'h0000;
            14'h0dbe: oData <= 16'h0000;
            14'h0dbf: oData <= 16'h0000;
            14'h0dc0: oData <= 16'h0000;
            14'h0dc1: oData <= 16'h0000;
            14'h0dc2: oData <= 16'h0000;
            14'h0dc3: oData <= 16'h0000;
            14'h0dc4: oData <= 16'h0000;
            14'h0dc5: oData <= 16'h2aa8;
            14'h0dc6: oData <= 16'hea00;
            14'h0dc7: oData <= 16'haffb;
            14'h0dc8: oData <= 16'hbfff;
            14'h0dc9: oData <= 16'hffaa;
            14'h0dca: oData <= 16'hffff;
            14'h0dcb: oData <= 16'hfffa;
            14'h0dcc: oData <= 16'hffaf;
            14'h0dcd: oData <= 16'hafeb;
            14'h0dce: oData <= 16'hebbf;
            14'h0dcf: oData <= 16'hafff;
            14'h0dd0: oData <= 16'h0000;
            14'h0dd1: oData <= 16'h0000;
            14'h0dd2: oData <= 16'h0000;
            14'h0dd3: oData <= 16'h0000;
            14'h0dd4: oData <= 16'h0000;
            14'h0dd5: oData <= 16'h0000;
            14'h0dd6: oData <= 16'h0000;
            14'h0dd7: oData <= 16'h0000;
            14'h0dd8: oData <= 16'h0000;
            14'h0dd9: oData <= 16'h2aa0;
            14'h0dda: oData <= 16'ha800;
            14'h0ddb: oData <= 16'hffaf;
            14'h0ddc: oData <= 16'hfffb;
            14'h0ddd: oData <= 16'heaab;
            14'h0dde: oData <= 16'hffff;
            14'h0ddf: oData <= 16'hfffa;
            14'h0de0: oData <= 16'hffaf;
            14'h0de1: oData <= 16'habea;
            14'h0de2: oData <= 16'heaff;
            14'h0de3: oData <= 16'hafff;
            14'h0de4: oData <= 16'h0000;
            14'h0de5: oData <= 16'h0000;
            14'h0de6: oData <= 16'h0000;
            14'h0de7: oData <= 16'h0000;
            14'h0de8: oData <= 16'h0000;
            14'h0de9: oData <= 16'h0000;
            14'h0dea: oData <= 16'h0000;
            14'h0deb: oData <= 16'h0000;
            14'h0dec: oData <= 16'h0000;
            14'h0ded: oData <= 16'haaa0;
            14'h0dee: oData <= 16'ha000;
            14'h0def: oData <= 16'hfafe;
            14'h0df0: oData <= 16'hffaf;
            14'h0df1: oData <= 16'haabf;
            14'h0df2: oData <= 16'hfffa;
            14'h0df3: oData <= 16'hfffa;
            14'h0df4: oData <= 16'hffab;
            14'h0df5: oData <= 16'haffa;
            14'h0df6: oData <= 16'hfeaa;
            14'h0df7: oData <= 16'hafff;
            14'h0df8: oData <= 16'h0000;
            14'h0df9: oData <= 16'h0000;
            14'h0dfa: oData <= 16'h0000;
            14'h0dfb: oData <= 16'h0000;
            14'h0dfc: oData <= 16'h0000;
            14'h0dfd: oData <= 16'h0000;
            14'h0dfe: oData <= 16'h0000;
            14'h0dff: oData <= 16'h0000;
            14'h0e00: oData <= 16'h0000;
            14'h0e01: oData <= 16'haa80;
            14'h0e02: oData <= 16'h8000;
            14'h0e03: oData <= 16'hafea;
            14'h0e04: oData <= 16'hfaff;
            14'h0e05: oData <= 16'hafff;
            14'h0e06: oData <= 16'haaaa;
            14'h0e07: oData <= 16'hffea;
            14'h0e08: oData <= 16'hbfeb;
            14'h0e09: oData <= 16'haaaa;
            14'h0e0a: oData <= 16'hffaa;
            14'h0e0b: oData <= 16'hafff;
            14'h0e0c: oData <= 16'h0000;
            14'h0e0d: oData <= 16'h0000;
            14'h0e0e: oData <= 16'h0000;
            14'h0e0f: oData <= 16'h0000;
            14'h0e10: oData <= 16'h0000;
            14'h0e11: oData <= 16'h0000;
            14'h0e12: oData <= 16'h0000;
            14'h0e13: oData <= 16'h0000;
            14'h0e14: oData <= 16'h0000;
            14'h0e15: oData <= 16'haa80;
            14'h0e16: oData <= 16'h0002;
            14'h0e17: oData <= 16'hffaa;
            14'h0e18: oData <= 16'haffa;
            14'h0e19: oData <= 16'hffff;
            14'h0e1a: oData <= 16'haaab;
            14'h0e1b: oData <= 16'haaaa;
            14'h0e1c: oData <= 16'haaaa;
            14'h0e1d: oData <= 16'haaaa;
            14'h0e1e: oData <= 16'hffff;
            14'h0e1f: oData <= 16'hafff;
            14'h0e20: oData <= 16'h0000;
            14'h0e21: oData <= 16'h0000;
            14'h0e22: oData <= 16'h0000;
            14'h0e23: oData <= 16'h0000;
            14'h0e24: oData <= 16'h0000;
            14'h0e25: oData <= 16'h0000;
            14'h0e26: oData <= 16'h0000;
            14'h0e27: oData <= 16'h0000;
            14'h0e28: oData <= 16'h0000;
            14'h0e29: oData <= 16'haa00;
            14'h0e2a: oData <= 16'h0002;
            14'h0e2b: oData <= 16'hfaa0;
            14'h0e2c: oData <= 16'hffaf;
            14'h0e2d: oData <= 16'hfffa;
            14'h0e2e: oData <= 16'hffff;
            14'h0e2f: oData <= 16'haaaf;
            14'h0e30: oData <= 16'haaaa;
            14'h0e31: oData <= 16'hffff;
            14'h0e32: oData <= 16'hffff;
            14'h0e33: oData <= 16'hafff;
            14'h0e34: oData <= 16'h0000;
            14'h0e35: oData <= 16'h0000;
            14'h0e36: oData <= 16'h0000;
            14'h0e37: oData <= 16'h0000;
            14'h0e38: oData <= 16'h0000;
            14'h0e39: oData <= 16'h0000;
            14'h0e3a: oData <= 16'h0000;
            14'h0e3b: oData <= 16'h0000;
            14'h0e3c: oData <= 16'h0000;
            14'h0e3d: oData <= 16'haa00;
            14'h0e3e: oData <= 16'h000a;
            14'h0e3f: oData <= 16'haa80;
            14'h0e40: oData <= 16'hfaff;
            14'h0e41: oData <= 16'hfeaf;
            14'h0e42: oData <= 16'hffff;
            14'h0e43: oData <= 16'hffff;
            14'h0e44: oData <= 16'hffff;
            14'h0e45: oData <= 16'hffff;
            14'h0e46: oData <= 16'hfbff;
            14'h0e47: oData <= 16'hafff;
            14'h0e48: oData <= 16'h0002;
            14'h0e49: oData <= 16'h0000;
            14'h0e4a: oData <= 16'h0000;
            14'h0e4b: oData <= 16'h0000;
            14'h0e4c: oData <= 16'h0000;
            14'h0e4d: oData <= 16'h0000;
            14'h0e4e: oData <= 16'h0000;
            14'h0e4f: oData <= 16'h0000;
            14'h0e50: oData <= 16'h0000;
            14'h0e51: oData <= 16'ha800;
            14'h0e52: oData <= 16'h000a;
            14'h0e53: oData <= 16'ha800;
            14'h0e54: oData <= 16'haffa;
            14'h0e55: oData <= 16'habff;
            14'h0e56: oData <= 16'hffff;
            14'h0e57: oData <= 16'hffff;
            14'h0e58: oData <= 16'hffff;
            14'h0e59: oData <= 16'hffff;
            14'h0e5a: oData <= 16'hfeff;
            14'h0e5b: oData <= 16'hbffb;
            14'h0e5c: oData <= 16'h0002;
            14'h0e5d: oData <= 16'h0000;
            14'h0e5e: oData <= 16'h0000;
            14'h0e5f: oData <= 16'h0000;
            14'h0e60: oData <= 16'h0000;
            14'h0e61: oData <= 16'h0000;
            14'h0e62: oData <= 16'h0000;
            14'h0e63: oData <= 16'h0000;
            14'h0e64: oData <= 16'h0000;
            14'h0e65: oData <= 16'ha800;
            14'h0e66: oData <= 16'h002a;
            14'h0e67: oData <= 16'h8000;
            14'h0e68: oData <= 16'hffaa;
            14'h0e69: oData <= 16'hffea;
            14'h0e6a: oData <= 16'hfffa;
            14'h0e6b: oData <= 16'haaaf;
            14'h0e6c: oData <= 16'haaaa;
            14'h0e6d: oData <= 16'hfffa;
            14'h0e6e: oData <= 16'hffaf;
            14'h0e6f: oData <= 16'hbffb;
            14'h0e70: oData <= 16'h0002;
            14'h0e71: oData <= 16'h0000;
            14'h0e72: oData <= 16'h0000;
            14'h0e73: oData <= 16'h0000;
            14'h0e74: oData <= 16'h0000;
            14'h0e75: oData <= 16'h0000;
            14'h0e76: oData <= 16'h0000;
            14'h0e77: oData <= 16'h0000;
            14'h0e78: oData <= 16'h0000;
            14'h0e79: oData <= 16'ha000;
            14'h0e7a: oData <= 16'h002a;
            14'h0e7b: oData <= 16'h0000;
            14'h0e7c: oData <= 16'hfaa8;
            14'h0e7d: oData <= 16'hfabf;
            14'h0e7e: oData <= 16'heaaf;
            14'h0e7f: oData <= 16'hffff;
            14'h0e80: oData <= 16'hffff;
            14'h0e81: oData <= 16'hffff;
            14'h0e82: oData <= 16'hfffb;
            14'h0e83: oData <= 16'hbffb;
            14'h0e84: oData <= 16'h0002;
            14'h0e85: oData <= 16'h0000;
            14'h0e86: oData <= 16'h0000;
            14'h0e87: oData <= 16'h0000;
            14'h0e88: oData <= 16'h0000;
            14'h0e89: oData <= 16'h0000;
            14'h0e8a: oData <= 16'h0000;
            14'h0e8b: oData <= 16'h0000;
            14'h0e8c: oData <= 16'h0000;
            14'h0e8d: oData <= 16'ha000;
            14'h0e8e: oData <= 16'h002a;
            14'h0e8f: oData <= 16'h0000;
            14'h0e90: oData <= 16'haa80;
            14'h0e91: oData <= 16'haffe;
            14'h0e92: oData <= 16'hbffe;
            14'h0e93: oData <= 16'haaaa;
            14'h0e94: oData <= 16'hfffa;
            14'h0e95: oData <= 16'habff;
            14'h0e96: oData <= 16'hfffe;
            14'h0e97: oData <= 16'hbffe;
            14'h0e98: oData <= 16'h0002;
            14'h0e99: oData <= 16'h0000;
            14'h0e9a: oData <= 16'h0000;
            14'h0e9b: oData <= 16'h0000;
            14'h0e9c: oData <= 16'h0000;
            14'h0e9d: oData <= 16'h0000;
            14'h0e9e: oData <= 16'h0000;
            14'h0e9f: oData <= 16'h0000;
            14'h0ea0: oData <= 16'h0000;
            14'h0ea1: oData <= 16'ha000;
            14'h0ea2: oData <= 16'h00aa;
            14'h0ea3: oData <= 16'h0000;
            14'h0ea4: oData <= 16'ha800;
            14'h0ea5: oData <= 16'hffea;
            14'h0ea6: oData <= 16'hfaab;
            14'h0ea7: oData <= 16'hffff;
            14'h0ea8: oData <= 16'haaaf;
            14'h0ea9: oData <= 16'hfeaa;
            14'h0eaa: oData <= 16'hafff;
            14'h0eab: oData <= 16'hbfff;
            14'h0eac: oData <= 16'h0002;
            14'h0ead: oData <= 16'h0000;
            14'h0eae: oData <= 16'h0000;
            14'h0eaf: oData <= 16'h0000;
            14'h0eb0: oData <= 16'h0000;
            14'h0eb1: oData <= 16'h0000;
            14'h0eb2: oData <= 16'h0000;
            14'h0eb3: oData <= 16'h0000;
            14'h0eb4: oData <= 16'h0000;
            14'h0eb5: oData <= 16'h8000;
            14'h0eb6: oData <= 16'h00aa;
            14'h0eb7: oData <= 16'h0000;
            14'h0eb8: oData <= 16'h0000;
            14'h0eb9: oData <= 16'hfeaa;
            14'h0eba: oData <= 16'hafff;
            14'h0ebb: oData <= 16'hffaa;
            14'h0ebc: oData <= 16'hffff;
            14'h0ebd: oData <= 16'hffff;
            14'h0ebe: oData <= 16'hfbff;
            14'h0ebf: oData <= 16'hbfff;
            14'h0ec0: oData <= 16'h0002;
            14'h0ec1: oData <= 16'h0000;
            14'h0ec2: oData <= 16'h0000;
            14'h0ec3: oData <= 16'h0000;
            14'h0ec4: oData <= 16'h0000;
            14'h0ec5: oData <= 16'h0000;
            14'h0ec6: oData <= 16'h0000;
            14'h0ec7: oData <= 16'h0000;
            14'h0ec8: oData <= 16'h0000;
            14'h0ec9: oData <= 16'h8000;
            14'h0eca: oData <= 16'h02aa;
            14'h0ecb: oData <= 16'h0000;
            14'h0ecc: oData <= 16'h0000;
            14'h0ecd: oData <= 16'heaa0;
            14'h0ece: oData <= 16'hffff;
            14'h0ecf: oData <= 16'haaff;
            14'h0ed0: oData <= 16'hfaaa;
            14'h0ed1: oData <= 16'hffff;
            14'h0ed2: oData <= 16'hfeab;
            14'h0ed3: oData <= 16'hafff;
            14'h0ed4: oData <= 16'h0002;
            14'h0ed5: oData <= 16'h0000;
            14'h0ed6: oData <= 16'h0000;
            14'h0ed7: oData <= 16'h0000;
            14'h0ed8: oData <= 16'h0000;
            14'h0ed9: oData <= 16'h0000;
            14'h0eda: oData <= 16'h0000;
            14'h0edb: oData <= 16'h0000;
            14'h0edc: oData <= 16'h0000;
            14'h0edd: oData <= 16'h0000;
            14'h0ede: oData <= 16'h02aa;
            14'h0edf: oData <= 16'h0000;
            14'h0ee0: oData <= 16'h0000;
            14'h0ee1: oData <= 16'haa00;
            14'h0ee2: oData <= 16'hfffa;
            14'h0ee3: oData <= 16'hffff;
            14'h0ee4: oData <= 16'hafff;
            14'h0ee5: oData <= 16'haaaa;
            14'h0ee6: oData <= 16'hfffe;
            14'h0ee7: oData <= 16'hafff;
            14'h0ee8: oData <= 16'h0a80;
            14'h0ee9: oData <= 16'h0000;
            14'h0eea: oData <= 16'h0000;
            14'h0eeb: oData <= 16'h0000;
            14'h0eec: oData <= 16'h0000;
            14'h0eed: oData <= 16'h0000;
            14'h0eee: oData <= 16'h0000;
            14'h0eef: oData <= 16'h0000;
            14'h0ef0: oData <= 16'h0000;
            14'h0ef1: oData <= 16'h0000;
            14'h0ef2: oData <= 16'h0aaa;
            14'h0ef3: oData <= 16'h0000;
            14'h0ef4: oData <= 16'h0000;
            14'h0ef5: oData <= 16'ha000;
            14'h0ef6: oData <= 16'hffea;
            14'h0ef7: oData <= 16'hffff;
            14'h0ef8: oData <= 16'hffff;
            14'h0ef9: oData <= 16'hffff;
            14'h0efa: oData <= 16'hffff;
            14'h0efb: oData <= 16'habff;
            14'h0efc: oData <= 16'h2aa0;
            14'h0efd: oData <= 16'h0000;
            14'h0efe: oData <= 16'h0000;
            14'h0eff: oData <= 16'h0000;
            14'h0f00: oData <= 16'h0000;
            14'h0f01: oData <= 16'h0000;
            14'h0f02: oData <= 16'h0000;
            14'h0f03: oData <= 16'h0000;
            14'h0f04: oData <= 16'h0000;
            14'h0f05: oData <= 16'h0000;
            14'h0f06: oData <= 16'h0aa8;
            14'h0f07: oData <= 16'h0000;
            14'h0f08: oData <= 16'h0000;
            14'h0f09: oData <= 16'ha000;
            14'h0f0a: oData <= 16'hfeaa;
            14'h0f0b: oData <= 16'hffff;
            14'h0f0c: oData <= 16'hffff;
            14'h0f0d: oData <= 16'hffff;
            14'h0f0e: oData <= 16'hffff;
            14'h0f0f: oData <= 16'h2bff;
            14'h0f10: oData <= 16'h2aa8;
            14'h0f11: oData <= 16'h0000;
            14'h0f12: oData <= 16'h0000;
            14'h0f13: oData <= 16'h0000;
            14'h0f14: oData <= 16'h0000;
            14'h0f15: oData <= 16'h0000;
            14'h0f16: oData <= 16'h0000;
            14'h0f17: oData <= 16'h0000;
            14'h0f18: oData <= 16'h0000;
            14'h0f19: oData <= 16'h0000;
            14'h0f1a: oData <= 16'h2aa8;
            14'h0f1b: oData <= 16'h0000;
            14'h0f1c: oData <= 16'h0000;
            14'h0f1d: oData <= 16'ha000;
            14'h0f1e: oData <= 16'haaaa;
            14'h0f1f: oData <= 16'hfffa;
            14'h0f20: oData <= 16'hffff;
            14'h0f21: oData <= 16'hffff;
            14'h0f22: oData <= 16'hffff;
            14'h0f23: oData <= 16'h2aff;
            14'h0f24: oData <= 16'h0aa8;
            14'h0f25: oData <= 16'h0000;
            14'h0f26: oData <= 16'h0000;
            14'h0f27: oData <= 16'h0000;
            14'h0f28: oData <= 16'h0000;
            14'h0f29: oData <= 16'h0000;
            14'h0f2a: oData <= 16'h0000;
            14'h0f2b: oData <= 16'h0000;
            14'h0f2c: oData <= 16'h0000;
            14'h0f2d: oData <= 16'h0000;
            14'h0f2e: oData <= 16'h2aa0;
            14'h0f2f: oData <= 16'h0000;
            14'h0f30: oData <= 16'h0000;
            14'h0f31: oData <= 16'ha000;
            14'h0f32: oData <= 16'haa2a;
            14'h0f33: oData <= 16'hfaaa;
            14'h0f34: oData <= 16'hffff;
            14'h0f35: oData <= 16'hffff;
            14'h0f36: oData <= 16'hffff;
            14'h0f37: oData <= 16'h0aaf;
            14'h0f38: oData <= 16'h02aa;
            14'h0f39: oData <= 16'h0000;
            14'h0f3a: oData <= 16'h0000;
            14'h0f3b: oData <= 16'h0000;
            14'h0f3c: oData <= 16'h0000;
            14'h0f3d: oData <= 16'h0000;
            14'h0f3e: oData <= 16'h0000;
            14'h0f3f: oData <= 16'h0000;
            14'h0f40: oData <= 16'h0000;
            14'h0f41: oData <= 16'h0000;
            14'h0f42: oData <= 16'haaa0;
            14'h0f43: oData <= 16'h0000;
            14'h0f44: oData <= 16'h0000;
            14'h0f45: oData <= 16'ha000;
            14'h0f46: oData <= 16'h002a;
            14'h0f47: oData <= 16'haaa8;
            14'h0f48: oData <= 16'hfffa;
            14'h0f49: oData <= 16'hffff;
            14'h0f4a: oData <= 16'hffff;
            14'h0f4b: oData <= 16'h82ab;
            14'h0f4c: oData <= 16'h02aa;
            14'h0f4d: oData <= 16'h0000;
            14'h0f4e: oData <= 16'h0000;
            14'h0f4f: oData <= 16'h0000;
            14'h0f50: oData <= 16'h0000;
            14'h0f51: oData <= 16'h0000;
            14'h0f52: oData <= 16'h0000;
            14'h0f53: oData <= 16'h0000;
            14'h0f54: oData <= 16'h0000;
            14'h0f55: oData <= 16'h0000;
            14'h0f56: oData <= 16'haa80;
            14'h0f57: oData <= 16'h0002;
            14'h0f58: oData <= 16'h0000;
            14'h0f59: oData <= 16'ha800;
            14'h0f5a: oData <= 16'h002a;
            14'h0f5b: oData <= 16'ha800;
            14'h0f5c: oData <= 16'hfaaa;
            14'h0f5d: oData <= 16'hffff;
            14'h0f5e: oData <= 16'hafff;
            14'h0f5f: oData <= 16'h802a;
            14'h0f60: oData <= 16'h00aa;
            14'h0f61: oData <= 16'h0000;
            14'h0f62: oData <= 16'h0000;
            14'h0f63: oData <= 16'h0000;
            14'h0f64: oData <= 16'h0000;
            14'h0f65: oData <= 16'h0000;
            14'h0f66: oData <= 16'h0000;
            14'h0f67: oData <= 16'h0000;
            14'h0f68: oData <= 16'h0000;
            14'h0f69: oData <= 16'h0000;
            14'h0f6a: oData <= 16'haa80;
            14'h0f6b: oData <= 16'h00aa;
            14'h0f6c: oData <= 16'h0000;
            14'h0f6d: oData <= 16'ha800;
            14'h0f6e: oData <= 16'h000a;
            14'h0f6f: oData <= 16'h0000;
            14'h0f70: oData <= 16'haaa8;
            14'h0f71: oData <= 16'haaaa;
            14'h0f72: oData <= 16'haaaa;
            14'h0f73: oData <= 16'ha002;
            14'h0f74: oData <= 16'h002a;
            14'h0f75: oData <= 16'h0000;
            14'h0f76: oData <= 16'h0000;
            14'h0f77: oData <= 16'h0000;
            14'h0f78: oData <= 16'h0000;
            14'h0f79: oData <= 16'h0000;
            14'h0f7a: oData <= 16'h0000;
            14'h0f7b: oData <= 16'h0000;
            14'h0f7c: oData <= 16'h0000;
            14'h0f7d: oData <= 16'h0000;
            14'h0f7e: oData <= 16'haa80;
            14'h0f7f: oData <= 16'h0aaa;
            14'h0f80: oData <= 16'h0000;
            14'h0f81: oData <= 16'ha800;
            14'h0f82: oData <= 16'h000a;
            14'h0f83: oData <= 16'h0000;
            14'h0f84: oData <= 16'ha800;
            14'h0f85: oData <= 16'haaaa;
            14'h0f86: oData <= 16'h2aaa;
            14'h0f87: oData <= 16'ha800;
            14'h0f88: oData <= 16'h002a;
            14'h0f89: oData <= 16'h0000;
            14'h0f8a: oData <= 16'h0000;
            14'h0f8b: oData <= 16'h0000;
            14'h0f8c: oData <= 16'h0000;
            14'h0f8d: oData <= 16'h0000;
            14'h0f8e: oData <= 16'h0000;
            14'h0f8f: oData <= 16'h0000;
            14'h0f90: oData <= 16'h0000;
            14'h0f91: oData <= 16'h0000;
            14'h0f92: oData <= 16'haa00;
            14'h0f93: oData <= 16'haaaa;
            14'h0f94: oData <= 16'h0002;
            14'h0f95: oData <= 16'ha800;
            14'h0f96: oData <= 16'h000a;
            14'h0f97: oData <= 16'h0000;
            14'h0f98: oData <= 16'h0000;
            14'h0f99: oData <= 16'h0000;
            14'h0f9a: oData <= 16'h0000;
            14'h0f9b: oData <= 16'haa00;
            14'h0f9c: oData <= 16'h000a;
            14'h0f9d: oData <= 16'h0000;
            14'h0f9e: oData <= 16'h0000;
            14'h0f9f: oData <= 16'h0000;
            14'h0fa0: oData <= 16'h0000;
            14'h0fa1: oData <= 16'h0000;
            14'h0fa2: oData <= 16'h0000;
            14'h0fa3: oData <= 16'h0000;
            14'h0fa4: oData <= 16'h0000;
            14'h0fa5: oData <= 16'h0000;
            14'h0fa6: oData <= 16'ha800;
            14'h0fa7: oData <= 16'haaaa;
            14'h0fa8: oData <= 16'h002a;
            14'h0fa9: oData <= 16'haa00;
            14'h0faa: oData <= 16'h000a;
            14'h0fab: oData <= 16'h0000;
            14'h0fac: oData <= 16'h0000;
            14'h0fad: oData <= 16'h0000;
            14'h0fae: oData <= 16'h0000;
            14'h0faf: oData <= 16'haaa0;
            14'h0fb0: oData <= 16'h0002;
            14'h0fb1: oData <= 16'h0000;
            14'h0fb2: oData <= 16'h0000;
            14'h0fb3: oData <= 16'h0000;
            14'h0fb4: oData <= 16'h0000;
            14'h0fb5: oData <= 16'h0000;
            14'h0fb6: oData <= 16'h0000;
            14'h0fb7: oData <= 16'h0000;
            14'h0fb8: oData <= 16'h0000;
            14'h0fb9: oData <= 16'h0000;
            14'h0fba: oData <= 16'h0000;
            14'h0fbb: oData <= 16'haaaa;
            14'h0fbc: oData <= 16'h0aaa;
            14'h0fbd: oData <= 16'haa00;
            14'h0fbe: oData <= 16'h0002;
            14'h0fbf: oData <= 16'h0000;
            14'h0fc0: oData <= 16'h0000;
            14'h0fc1: oData <= 16'h0000;
            14'h0fc2: oData <= 16'h0000;
            14'h0fc3: oData <= 16'haaa8;
            14'h0fc4: oData <= 16'h000a;
            14'h0fc5: oData <= 16'h0000;
            14'h0fc6: oData <= 16'h0000;
            14'h0fc7: oData <= 16'h0000;
            14'h0fc8: oData <= 16'h0000;
            14'h0fc9: oData <= 16'h0000;
            14'h0fca: oData <= 16'h0000;
            14'h0fcb: oData <= 16'h0000;
            14'h0fcc: oData <= 16'h0000;
            14'h0fcd: oData <= 16'h0000;
            14'h0fce: oData <= 16'h0000;
            14'h0fcf: oData <= 16'haa80;
            14'h0fd0: oData <= 16'haaaa;
            14'h0fd1: oData <= 16'haa00;
            14'h0fd2: oData <= 16'h0002;
            14'h0fd3: oData <= 16'h0000;
            14'h0fd4: oData <= 16'h0000;
            14'h0fd5: oData <= 16'h0000;
            14'h0fd6: oData <= 16'h0000;
            14'h0fd7: oData <= 16'haaaa;
            14'h0fd8: oData <= 16'h000a;
            14'h0fd9: oData <= 16'h0000;
            14'h0fda: oData <= 16'h0000;
            14'h0fdb: oData <= 16'h0000;
            14'h0fdc: oData <= 16'h0000;
            14'h0fdd: oData <= 16'h0000;
            14'h0fde: oData <= 16'h0000;
            14'h0fdf: oData <= 16'h0000;
            14'h0fe0: oData <= 16'h0000;
            14'h0fe1: oData <= 16'h0000;
            14'h0fe2: oData <= 16'h0000;
            14'h0fe3: oData <= 16'ha800;
            14'h0fe4: oData <= 16'haaaa;
            14'h0fe5: oData <= 16'haa2a;
            14'h0fe6: oData <= 16'h0002;
            14'h0fe7: oData <= 16'h0000;
            14'h0fe8: oData <= 16'h0000;
            14'h0fe9: oData <= 16'h0000;
            14'h0fea: oData <= 16'ha800;
            14'h0feb: oData <= 16'haaaa;
            14'h0fec: oData <= 16'h000a;
            14'h0fed: oData <= 16'h0000;
            14'h0fee: oData <= 16'h0000;
            14'h0fef: oData <= 16'h0000;
            14'h0ff0: oData <= 16'h0000;
            14'h0ff1: oData <= 16'h0000;
            14'h0ff2: oData <= 16'h0000;
            14'h0ff3: oData <= 16'h0000;
            14'h0ff4: oData <= 16'h0000;
            14'h0ff5: oData <= 16'h0000;
            14'h0ff6: oData <= 16'h0000;
            14'h0ff7: oData <= 16'h0000;
            14'h0ff8: oData <= 16'haaaa;
            14'h0ff9: oData <= 16'haaaa;
            14'h0ffa: oData <= 16'h0002;
            14'h0ffb: oData <= 16'h0000;
            14'h0ffc: oData <= 16'h0000;
            14'h0ffd: oData <= 16'h0000;
            14'h0ffe: oData <= 16'haaa8;
            14'h0fff: oData <= 16'haaaa;
            14'h1000: oData <= 16'h0002;
            14'h1001: oData <= 16'h0000;
            14'h1002: oData <= 16'h0000;
            14'h1003: oData <= 16'h0000;
            14'h1004: oData <= 16'h0000;
            14'h1005: oData <= 16'h0000;
            14'h1006: oData <= 16'h0000;
            14'h1007: oData <= 16'h0000;
            14'h1008: oData <= 16'h0000;
            14'h1009: oData <= 16'h0000;
            14'h100a: oData <= 16'h0000;
            14'h100b: oData <= 16'h0000;
            14'h100c: oData <= 16'haaa0;
            14'h100d: oData <= 16'haaaa;
            14'h100e: oData <= 16'h2aaa;
            14'h100f: oData <= 16'h0000;
            14'h1010: oData <= 16'h0000;
            14'h1011: oData <= 16'ha000;
            14'h1012: oData <= 16'haaaa;
            14'h1013: oData <= 16'haaaa;
            14'h1014: oData <= 16'h0000;
            14'h1015: oData <= 16'h0000;
            14'h1016: oData <= 16'h0000;
            14'h1017: oData <= 16'h0000;
            14'h1018: oData <= 16'h0000;
            14'h1019: oData <= 16'h0000;
            14'h101a: oData <= 16'h0000;
            14'h101b: oData <= 16'h0000;
            14'h101c: oData <= 16'h0000;
            14'h101d: oData <= 16'h0000;
            14'h101e: oData <= 16'h0000;
            14'h101f: oData <= 16'h0000;
            14'h1020: oData <= 16'ha800;
            14'h1021: oData <= 16'haaaa;
            14'h1022: oData <= 16'haaaa;
            14'h1023: oData <= 16'h2aaa;
            14'h1024: oData <= 16'h0000;
            14'h1025: oData <= 16'haaa0;
            14'h1026: oData <= 16'haaaa;
            14'h1027: oData <= 16'haaaa;
            14'h1028: oData <= 16'h0000;
            14'h1029: oData <= 16'ha000;
            14'h102a: oData <= 16'h00aa;
            14'h102b: oData <= 16'h0000;
            14'h102c: oData <= 16'h0000;
            14'h102d: oData <= 16'h0000;
            14'h102e: oData <= 16'h0000;
            14'h102f: oData <= 16'h0000;
            14'h1030: oData <= 16'h0000;
            14'h1031: oData <= 16'h00a8;
            14'h1032: oData <= 16'h0000;
            14'h1033: oData <= 16'h0000;
            14'h1034: oData <= 16'h8000;
            14'h1035: oData <= 16'haaaa;
            14'h1036: oData <= 16'haaaa;
            14'h1037: oData <= 16'haaaa;
            14'h1038: oData <= 16'haaaa;
            14'h1039: oData <= 16'haaaa;
            14'h103a: oData <= 16'haaaa;
            14'h103b: oData <= 16'haa82;
            14'h103c: oData <= 16'h0002;
            14'h103d: oData <= 16'haa80;
            14'h103e: oData <= 16'h02aa;
            14'h103f: oData <= 16'h0000;
            14'h1040: oData <= 16'h0000;
            14'h1041: oData <= 16'h0000;
            14'h1042: oData <= 16'h0000;
            14'h1043: oData <= 16'h0000;
            14'h1044: oData <= 16'h0000;
            14'h1045: oData <= 16'h02aa;
            14'h1046: oData <= 16'h0000;
            14'h1047: oData <= 16'h0000;
            14'h1048: oData <= 16'h0000;
            14'h1049: oData <= 16'haaa0;
            14'h104a: oData <= 16'haaaa;
            14'h104b: oData <= 16'haaaa;
            14'h104c: oData <= 16'haaaa;
            14'h104d: oData <= 16'haaaa;
            14'h104e: oData <= 16'h0aaa;
            14'h104f: oData <= 16'haa00;
            14'h1050: oData <= 16'h000a;
            14'h1051: oData <= 16'haaa0;
            14'h1052: oData <= 16'h0aaa;
            14'h1053: oData <= 16'h0000;
            14'h1054: oData <= 16'h0000;
            14'h1055: oData <= 16'h0000;
            14'h1056: oData <= 16'h0000;
            14'h1057: oData <= 16'h0000;
            14'h1058: oData <= 16'h0000;
            14'h1059: oData <= 16'h02aa;
            14'h105a: oData <= 16'h0000;
            14'h105b: oData <= 16'h0000;
            14'h105c: oData <= 16'h0000;
            14'h105d: oData <= 16'haaa0;
            14'h105e: oData <= 16'haaaa;
            14'h105f: oData <= 16'haaaa;
            14'h1060: oData <= 16'haaaa;
            14'h1061: oData <= 16'haaaa;
            14'h1062: oData <= 16'h000a;
            14'h1063: oData <= 16'ha800;
            14'h1064: oData <= 16'h002a;
            14'h1065: oData <= 16'haaa8;
            14'h1066: oData <= 16'h2aaa;
            14'h1067: oData <= 16'h0000;
            14'h1068: oData <= 16'h0000;
            14'h1069: oData <= 16'h0000;
            14'h106a: oData <= 16'h0000;
            14'h106b: oData <= 16'h0000;
            14'h106c: oData <= 16'h0000;
            14'h106d: oData <= 16'h0aaa;
            14'h106e: oData <= 16'h0000;
            14'h106f: oData <= 16'h0000;
            14'h1070: oData <= 16'h0000;
            14'h1071: oData <= 16'h2aa0;
            14'h1072: oData <= 16'ha000;
            14'h1073: oData <= 16'haaaa;
            14'h1074: oData <= 16'haaaa;
            14'h1075: oData <= 16'h2aaa;
            14'h1076: oData <= 16'h0000;
            14'h1077: oData <= 16'ha000;
            14'h1078: oData <= 16'h00aa;
            14'h1079: oData <= 16'h2aa8;
            14'h107a: oData <= 16'h2aa0;
            14'h107b: oData <= 16'h0000;
            14'h107c: oData <= 16'h0000;
            14'h107d: oData <= 16'h0000;
            14'h107e: oData <= 16'h0000;
            14'h107f: oData <= 16'h0000;
            14'h1080: oData <= 16'h0000;
            14'h1081: oData <= 16'h2aa8;
            14'h1082: oData <= 16'h0000;
            14'h1083: oData <= 16'h0000;
            14'h1084: oData <= 16'h0000;
            14'h1085: oData <= 16'h2aa0;
            14'h1086: oData <= 16'h0000;
            14'h1087: oData <= 16'ha000;
            14'h1088: oData <= 16'haaaa;
            14'h1089: oData <= 16'h002a;
            14'h108a: oData <= 16'h0000;
            14'h108b: oData <= 16'h8000;
            14'h108c: oData <= 16'h00aa;
            14'h108d: oData <= 16'h02aa;
            14'h108e: oData <= 16'h2aa0;
            14'h108f: oData <= 16'h0000;
            14'h1090: oData <= 16'h0000;
            14'h1091: oData <= 16'h0000;
            14'h1092: oData <= 16'h0000;
            14'h1093: oData <= 16'h0000;
            14'h1094: oData <= 16'h0000;
            14'h1095: oData <= 16'haaa0;
            14'h1096: oData <= 16'h0000;
            14'h1097: oData <= 16'h0000;
            14'h1098: oData <= 16'h0000;
            14'h1099: oData <= 16'h2aa8;
            14'h109a: oData <= 16'h0000;
            14'h109b: oData <= 16'h0000;
            14'h109c: oData <= 16'h0000;
            14'h109d: oData <= 16'h0000;
            14'h109e: oData <= 16'h0000;
            14'h109f: oData <= 16'h0000;
            14'h10a0: oData <= 16'h00aa;
            14'h10a1: oData <= 16'h02aa;
            14'h10a2: oData <= 16'h2aa0;
            14'h10a3: oData <= 16'h0000;
            14'h10a4: oData <= 16'h0000;
            14'h10a5: oData <= 16'h0000;
            14'h10a6: oData <= 16'h0000;
            14'h10a7: oData <= 16'h0000;
            14'h10a8: oData <= 16'h0000;
            14'h10a9: oData <= 16'haa80;
            14'h10aa: oData <= 16'h0000;
            14'h10ab: oData <= 16'h0000;
            14'h10ac: oData <= 16'h0000;
            14'h10ad: oData <= 16'h0aa8;
            14'h10ae: oData <= 16'h0000;
            14'h10af: oData <= 16'h0000;
            14'h10b0: oData <= 16'h0000;
            14'h10b1: oData <= 16'h0000;
            14'h10b2: oData <= 16'h0000;
            14'h10b3: oData <= 16'h0000;
            14'h10b4: oData <= 16'h0028;
            14'h10b5: oData <= 16'h00aa;
            14'h10b6: oData <= 16'h0aa8;
            14'h10b7: oData <= 16'h0000;
            14'h10b8: oData <= 16'h0000;
            14'h10b9: oData <= 16'h0000;
            14'h10ba: oData <= 16'h0000;
            14'h10bb: oData <= 16'h0000;
            14'h10bc: oData <= 16'h0000;
            14'h10bd: oData <= 16'haa80;
            14'h10be: oData <= 16'h0002;
            14'h10bf: oData <= 16'h0000;
            14'h10c0: oData <= 16'h0000;
            14'h10c1: oData <= 16'h0aa8;
            14'h10c2: oData <= 16'h0000;
            14'h10c3: oData <= 16'h00a8;
            14'h10c4: oData <= 16'h0000;
            14'h10c5: oData <= 16'h0000;
            14'h10c6: oData <= 16'h0000;
            14'h10c7: oData <= 16'h0000;
            14'h10c8: oData <= 16'h0000;
            14'h10c9: oData <= 16'h00aa;
            14'h10ca: oData <= 16'h0aa8;
            14'h10cb: oData <= 16'h0280;
            14'h10cc: oData <= 16'h0000;
            14'h10cd: oData <= 16'h0000;
            14'h10ce: oData <= 16'h0000;
            14'h10cf: oData <= 16'h0000;
            14'h10d0: oData <= 16'h0000;
            14'h10d1: oData <= 16'haa00;
            14'h10d2: oData <= 16'h000a;
            14'h10d3: oData <= 16'h0000;
            14'h10d4: oData <= 16'h0000;
            14'h10d5: oData <= 16'h0aa8;
            14'h10d6: oData <= 16'h0000;
            14'h10d7: oData <= 16'h02aa;
            14'h10d8: oData <= 16'h0000;
            14'h10d9: oData <= 16'h0000;
            14'h10da: oData <= 16'h0000;
            14'h10db: oData <= 16'h0000;
            14'h10dc: oData <= 16'h0000;
            14'h10dd: oData <= 16'ha0aa;
            14'h10de: oData <= 16'h02aa;
            14'h10df: oData <= 16'h0aa0;
            14'h10e0: oData <= 16'h0000;
            14'h10e1: oData <= 16'h0000;
            14'h10e2: oData <= 16'h0000;
            14'h10e3: oData <= 16'h0000;
            14'h10e4: oData <= 16'h0000;
            14'h10e5: oData <= 16'ha800;
            14'h10e6: oData <= 16'h000a;
            14'h10e7: oData <= 16'h0000;
            14'h10e8: oData <= 16'h0000;
            14'h10e9: oData <= 16'h0aaa;
            14'h10ea: oData <= 16'ha000;
            14'h10eb: oData <= 16'h02aa;
            14'h10ec: oData <= 16'h0000;
            14'h10ed: oData <= 16'h0000;
            14'h10ee: oData <= 16'h0000;
            14'h10ef: oData <= 16'h0000;
            14'h10f0: oData <= 16'h0000;
            14'h10f1: oData <= 16'haaaa;
            14'h10f2: oData <= 16'h02aa;
            14'h10f3: oData <= 16'h0aa0;
            14'h10f4: oData <= 16'h0000;
            14'h10f5: oData <= 16'h0000;
            14'h10f6: oData <= 16'h0000;
            14'h10f7: oData <= 16'h0000;
            14'h10f8: oData <= 16'h0000;
            14'h10f9: oData <= 16'ha800;
            14'h10fa: oData <= 16'h002a;
            14'h10fb: oData <= 16'h0000;
            14'h10fc: oData <= 16'h0000;
            14'h10fd: oData <= 16'h02aa;
            14'h10fe: oData <= 16'haa80;
            14'h10ff: oData <= 16'h0aaa;
            14'h1100: oData <= 16'h0000;
            14'h1101: oData <= 16'h0000;
            14'h1102: oData <= 16'h0000;
            14'h1103: oData <= 16'h0000;
            14'h1104: oData <= 16'h0000;
            14'h1105: oData <= 16'haaaa;
            14'h1106: oData <= 16'h00aa;
            14'h1107: oData <= 16'h0aa8;
            14'h1108: oData <= 16'h0000;
            14'h1109: oData <= 16'h0000;
            14'h110a: oData <= 16'h0000;
            14'h110b: oData <= 16'h0000;
            14'h110c: oData <= 16'h0000;
            14'h110d: oData <= 16'ha000;
            14'h110e: oData <= 16'h00aa;
            14'h110f: oData <= 16'h0000;
            14'h1110: oData <= 16'h0000;
            14'h1111: oData <= 16'h02aa;
            14'h1112: oData <= 16'haaa8;
            14'h1113: oData <= 16'h2aaa;
            14'h1114: oData <= 16'h0000;
            14'h1115: oData <= 16'h0000;
            14'h1116: oData <= 16'h0000;
            14'h1117: oData <= 16'h0000;
            14'h1118: oData <= 16'h0000;
            14'h1119: oData <= 16'haaa8;
            14'h111a: oData <= 16'h000a;
            14'h111b: oData <= 16'h0aa8;
            14'h111c: oData <= 16'h0000;
            14'h111d: oData <= 16'h0000;
            14'h111e: oData <= 16'h0000;
            14'h111f: oData <= 16'h0000;
            14'h1120: oData <= 16'h0000;
            14'h1121: oData <= 16'h8000;
            14'h1122: oData <= 16'h00aa;
            14'h1123: oData <= 16'h0000;
            14'h1124: oData <= 16'h0000;
            14'h1125: oData <= 16'ha2aa;
            14'h1126: oData <= 16'haaaa;
            14'h1127: oData <= 16'haaaa;
            14'h1128: oData <= 16'h0000;
            14'h1129: oData <= 16'h0000;
            14'h112a: oData <= 16'h0000;
            14'h112b: oData <= 16'h0000;
            14'h112c: oData <= 16'h0000;
            14'h112d: oData <= 16'haaa0;
            14'h112e: oData <= 16'h0000;
            14'h112f: oData <= 16'h02aa;
            14'h1130: oData <= 16'h0000;
            14'h1131: oData <= 16'h0000;
            14'h1132: oData <= 16'h0000;
            14'h1133: oData <= 16'h0000;
            14'h1134: oData <= 16'h0000;
            14'h1135: oData <= 16'h8000;
            14'h1136: oData <= 16'h02aa;
            14'h1137: oData <= 16'h0000;
            14'h1138: oData <= 16'h8000;
            14'h1139: oData <= 16'haaaa;
            14'h113a: oData <= 16'haaaa;
            14'h113b: oData <= 16'haa82;
            14'h113c: oData <= 16'h0002;
            14'h113d: oData <= 16'h0000;
            14'h113e: oData <= 16'h0000;
            14'h113f: oData <= 16'h0000;
            14'h1140: oData <= 16'h0000;
            14'h1141: oData <= 16'h0000;
            14'h1142: oData <= 16'h8000;
            14'h1143: oData <= 16'h02aa;
            14'h1144: oData <= 16'h0000;
            14'h1145: oData <= 16'h0000;
            14'h1146: oData <= 16'h0000;
            14'h1147: oData <= 16'h0000;
            14'h1148: oData <= 16'h0000;
            14'h1149: oData <= 16'h0000;
            14'h114a: oData <= 16'h0aaa;
            14'h114b: oData <= 16'h0000;
            14'h114c: oData <= 16'h8000;
            14'h114d: oData <= 16'haaaa;
            14'h114e: oData <= 16'h2aaa;
            14'h114f: oData <= 16'haa00;
            14'h1150: oData <= 16'h0002;
            14'h1151: oData <= 16'h0000;
            14'h1152: oData <= 16'h0000;
            14'h1153: oData <= 16'h0000;
            14'h1154: oData <= 16'h0000;
            14'h1155: oData <= 16'h0000;
            14'h1156: oData <= 16'ha000;
            14'h1157: oData <= 16'h00aa;
            14'h1158: oData <= 16'h0000;
            14'h1159: oData <= 16'h0000;
            14'h115a: oData <= 16'h0000;
            14'h115b: oData <= 16'h0000;
            14'h115c: oData <= 16'h0000;
            14'h115d: oData <= 16'h0000;
            14'h115e: oData <= 16'h0aa8;
            14'h115f: oData <= 16'h0000;
            14'h1160: oData <= 16'ha000;
            14'h1161: oData <= 16'haaaa;
            14'h1162: oData <= 16'h00aa;
            14'h1163: oData <= 16'haa00;
            14'h1164: oData <= 16'h000a;
            14'h1165: oData <= 16'h0000;
            14'h1166: oData <= 16'h0000;
            14'h1167: oData <= 16'h0000;
            14'h1168: oData <= 16'h0000;
            14'h1169: oData <= 16'h0000;
            14'h116a: oData <= 16'haa80;
            14'h116b: oData <= 16'h002a;
            14'h116c: oData <= 16'h0000;
            14'h116d: oData <= 16'h0000;
            14'h116e: oData <= 16'h0000;
            14'h116f: oData <= 16'h0000;
            14'h1170: oData <= 16'h0000;
            14'h1171: oData <= 16'h0000;
            14'h1172: oData <= 16'h2aa8;
            14'h1173: oData <= 16'h0000;
            14'h1174: oData <= 16'ha000;
            14'h1175: oData <= 16'haaaa;
            14'h1176: oData <= 16'h000a;
            14'h1177: oData <= 16'ha800;
            14'h1178: oData <= 16'h002a;
            14'h1179: oData <= 16'h0000;
            14'h117a: oData <= 16'h0000;
            14'h117b: oData <= 16'h0000;
            14'h117c: oData <= 16'h0000;
            14'h117d: oData <= 16'h0000;
            14'h117e: oData <= 16'haaaa;
            14'h117f: oData <= 16'h000a;
            14'h1180: oData <= 16'h0000;
            14'h1181: oData <= 16'h0000;
            14'h1182: oData <= 16'h0000;
            14'h1183: oData <= 16'h0000;
            14'h1184: oData <= 16'h0000;
            14'h1185: oData <= 16'h0000;
            14'h1186: oData <= 16'haaa0;
            14'h1187: oData <= 16'h0000;
            14'h1188: oData <= 16'ha800;
            14'h1189: oData <= 16'h2aaa;
            14'h118a: oData <= 16'h0000;
            14'h118b: oData <= 16'ha000;
            14'h118c: oData <= 16'h00aa;
            14'h118d: oData <= 16'h0000;
            14'h118e: oData <= 16'h0000;
            14'h118f: oData <= 16'h0000;
            14'h1190: oData <= 16'h0000;
            14'h1191: oData <= 16'h8000;
            14'h1192: oData <= 16'haaaa;
            14'h1193: oData <= 16'h0002;
            14'h1194: oData <= 16'h0000;
            14'h1195: oData <= 16'h0000;
            14'h1196: oData <= 16'h0000;
            14'h1197: oData <= 16'h0000;
            14'h1198: oData <= 16'h0000;
            14'h1199: oData <= 16'h0000;
            14'h119a: oData <= 16'haa80;
            14'h119b: oData <= 16'h0000;
            14'h119c: oData <= 16'haa00;
            14'h119d: oData <= 16'h02aa;
            14'h119e: oData <= 16'h0000;
            14'h119f: oData <= 16'h8000;
            14'h11a0: oData <= 16'h00aa;
            14'h11a1: oData <= 16'h0000;
            14'h11a2: oData <= 16'h0000;
            14'h11a3: oData <= 16'h0000;
            14'h11a4: oData <= 16'h0000;
            14'h11a5: oData <= 16'h8000;
            14'h11a6: oData <= 16'h2aaa;
            14'h11a7: oData <= 16'h0000;
            14'h11a8: oData <= 16'h0000;
            14'h11a9: oData <= 16'h0000;
            14'h11aa: oData <= 16'h0000;
            14'h11ab: oData <= 16'h0000;
            14'h11ac: oData <= 16'h0000;
            14'h11ad: oData <= 16'h0000;
            14'h11ae: oData <= 16'haa80;
            14'h11af: oData <= 16'h0002;
            14'h11b0: oData <= 16'haa80;
            14'h11b1: oData <= 16'h0002;
            14'h11b2: oData <= 16'h0000;
            14'h11b3: oData <= 16'h8000;
            14'h11b4: oData <= 16'h02aa;
            14'h11b5: oData <= 16'h0000;
            14'h11b6: oData <= 16'h0000;
            14'h11b7: oData <= 16'h0000;
            14'h11b8: oData <= 16'h0000;
            14'h11b9: oData <= 16'ha000;
            14'h11ba: oData <= 16'h02aa;
            14'h11bb: oData <= 16'h0000;
            14'h11bc: oData <= 16'h0000;
            14'h11bd: oData <= 16'h0000;
            14'h11be: oData <= 16'h0000;
            14'h11bf: oData <= 16'h0000;
            14'h11c0: oData <= 16'h0000;
            14'h11c1: oData <= 16'h0000;
            14'h11c2: oData <= 16'haa00;
            14'h11c3: oData <= 16'h000a;
            14'h11c4: oData <= 16'haaa8;
            14'h11c5: oData <= 16'h0000;
            14'h11c6: oData <= 16'h0000;
            14'h11c7: oData <= 16'h0000;
            14'h11c8: oData <= 16'h0aaa;
            14'h11c9: oData <= 16'h0000;
            14'h11ca: oData <= 16'h0000;
            14'h11cb: oData <= 16'h0000;
            14'h11cc: oData <= 16'h0000;
            14'h11cd: oData <= 16'ha000;
            14'h11ce: oData <= 16'h002a;
            14'h11cf: oData <= 16'h0000;
            14'h11d0: oData <= 16'h0000;
            14'h11d1: oData <= 16'h0000;
            14'h11d2: oData <= 16'h0000;
            14'h11d3: oData <= 16'h0000;
            14'h11d4: oData <= 16'h0000;
            14'h11d5: oData <= 16'h0000;
            14'h11d6: oData <= 16'ha800;
            14'h11d7: oData <= 16'h000a;
            14'h11d8: oData <= 16'h2aaa;
            14'h11d9: oData <= 16'h0000;
            14'h11da: oData <= 16'h0000;
            14'h11db: oData <= 16'h0000;
            14'h11dc: oData <= 16'h2aa8;
            14'h11dd: oData <= 16'h0000;
            14'h11de: oData <= 16'h0000;
            14'h11df: oData <= 16'h0000;
            14'h11e0: oData <= 16'h0000;
            14'h11e1: oData <= 16'ha000;
            14'h11e2: oData <= 16'h002a;
            14'h11e3: oData <= 16'h0000;
            14'h11e4: oData <= 16'h0000;
            14'h11e5: oData <= 16'h0000;
            14'h11e6: oData <= 16'h0000;
            14'h11e7: oData <= 16'h0000;
            14'h11e8: oData <= 16'h0000;
            14'h11e9: oData <= 16'h0000;
            14'h11ea: oData <= 16'ha800;
            14'h11eb: oData <= 16'h802a;
            14'h11ec: oData <= 16'h0aaa;
            14'h11ed: oData <= 16'h0000;
            14'h11ee: oData <= 16'h0000;
            14'h11ef: oData <= 16'h0000;
            14'h11f0: oData <= 16'h2aa0;
            14'h11f1: oData <= 16'h0000;
            14'h11f2: oData <= 16'h0000;
            14'h11f3: oData <= 16'h0000;
            14'h11f4: oData <= 16'h0000;
            14'h11f5: oData <= 16'ha000;
            14'h11f6: oData <= 16'h002a;
            14'h11f7: oData <= 16'h0000;
            14'h11f8: oData <= 16'h0000;
            14'h11f9: oData <= 16'h0000;
            14'h11fa: oData <= 16'h0000;
            14'h11fb: oData <= 16'h0000;
            14'h11fc: oData <= 16'h0000;
            14'h11fd: oData <= 16'h0000;
            14'h11fe: oData <= 16'ha000;
            14'h11ff: oData <= 16'ha0aa;
            14'h1200: oData <= 16'h02aa;
            14'h1201: oData <= 16'h0000;
            14'h1202: oData <= 16'h0000;
            14'h1203: oData <= 16'h0000;
            14'h1204: oData <= 16'haaa0;
            14'h1205: oData <= 16'h0000;
            14'h1206: oData <= 16'h0000;
            14'h1207: oData <= 16'h0000;
            14'h1208: oData <= 16'h0000;
            14'h1209: oData <= 16'h8000;
            14'h120a: oData <= 16'h00aa;
            14'h120b: oData <= 16'h0000;
            14'h120c: oData <= 16'h0000;
            14'h120d: oData <= 16'h0000;
            14'h120e: oData <= 16'h0000;
            14'h120f: oData <= 16'h0000;
            14'h1210: oData <= 16'h0000;
            14'h1211: oData <= 16'h0000;
            14'h1212: oData <= 16'h8000;
            14'h1213: oData <= 16'ha8aa;
            14'h1214: oData <= 16'h00aa;
            14'h1215: oData <= 16'h0000;
            14'h1216: oData <= 16'h0000;
            14'h1217: oData <= 16'h0000;
            14'h1218: oData <= 16'haa80;
            14'h1219: oData <= 16'h0002;
            14'h121a: oData <= 16'h0000;
            14'h121b: oData <= 16'h0000;
            14'h121c: oData <= 16'h0000;
            14'h121d: oData <= 16'h8000;
            14'h121e: oData <= 16'h02aa;
            14'h121f: oData <= 16'h0000;
            14'h1220: oData <= 16'h0000;
            14'h1221: oData <= 16'h0000;
            14'h1222: oData <= 16'h0000;
            14'h1223: oData <= 16'h0000;
            14'h1224: oData <= 16'h0000;
            14'h1225: oData <= 16'h0000;
            14'h1226: oData <= 16'h8000;
            14'h1227: oData <= 16'haaaa;
            14'h1228: oData <= 16'h000a;
            14'h1229: oData <= 16'h0000;
            14'h122a: oData <= 16'h0000;
            14'h122b: oData <= 16'h0000;
            14'h122c: oData <= 16'haa00;
            14'h122d: oData <= 16'h000a;
            14'h122e: oData <= 16'h0000;
            14'h122f: oData <= 16'h0000;
            14'h1230: oData <= 16'h0000;
            14'h1231: oData <= 16'h0000;
            14'h1232: oData <= 16'h02aa;
            14'h1233: oData <= 16'h0000;
            14'h1234: oData <= 16'h0000;
            14'h1235: oData <= 16'h0000;
            14'h1236: oData <= 16'h0000;
            14'h1237: oData <= 16'h0000;
            14'h1238: oData <= 16'h0000;
            14'h1239: oData <= 16'h0000;
            14'h123a: oData <= 16'h0000;
            14'h123b: oData <= 16'haaaa;
            14'h123c: oData <= 16'h0002;
            14'h123d: oData <= 16'h0000;
            14'h123e: oData <= 16'h0000;
            14'h123f: oData <= 16'h0000;
            14'h1240: oData <= 16'ha800;
            14'h1241: oData <= 16'h000a;
            14'h1242: oData <= 16'h0000;
            14'h1243: oData <= 16'h0000;
            14'h1244: oData <= 16'h0000;
            14'h1245: oData <= 16'h0000;
            14'h1246: oData <= 16'h0aa8;
            14'h1247: oData <= 16'h0000;
            14'h1248: oData <= 16'h0000;
            14'h1249: oData <= 16'h0000;
            14'h124a: oData <= 16'h0000;
            14'h124b: oData <= 16'h0000;
            14'h124c: oData <= 16'h0000;
            14'h124d: oData <= 16'h0000;
            14'h124e: oData <= 16'h0000;
            14'h124f: oData <= 16'haaa8;
            14'h1250: oData <= 16'h0000;
            14'h1251: oData <= 16'h0000;
            14'h1252: oData <= 16'h0000;
            14'h1253: oData <= 16'h0000;
            14'h1254: oData <= 16'ha800;
            14'h1255: oData <= 16'h002a;
            14'h1256: oData <= 16'h0000;
            14'h1257: oData <= 16'h0000;
            14'h1258: oData <= 16'h0000;
            14'h1259: oData <= 16'h0000;
            14'h125a: oData <= 16'h2aa8;
            14'h125b: oData <= 16'h0000;
            14'h125c: oData <= 16'h0000;
            14'h125d: oData <= 16'h0000;
            14'h125e: oData <= 16'h0000;
            14'h125f: oData <= 16'h0000;
            14'h1260: oData <= 16'h0000;
            14'h1261: oData <= 16'h0000;
            14'h1262: oData <= 16'h0000;
            14'h1263: oData <= 16'h2aa8;
            14'h1264: oData <= 16'h0000;
            14'h1265: oData <= 16'h0000;
            14'h1266: oData <= 16'h0000;
            14'h1267: oData <= 16'h0000;
            14'h1268: oData <= 16'ha000;
            14'h1269: oData <= 16'h00aa;
            14'h126a: oData <= 16'h0000;
            14'h126b: oData <= 16'h0000;
            14'h126c: oData <= 16'h0000;
            14'h126d: oData <= 16'h0000;
            14'h126e: oData <= 16'h2aa0;
            14'h126f: oData <= 16'h0000;
            14'h1270: oData <= 16'h0000;
            14'h1271: oData <= 16'h0000;
            14'h1272: oData <= 16'h0000;
            14'h1273: oData <= 16'h0000;
            14'h1274: oData <= 16'h0000;
            14'h1275: oData <= 16'h0000;
            14'h1276: oData <= 16'h0000;
            14'h1277: oData <= 16'h0aa0;
            14'h1278: oData <= 16'h0000;
            14'h1279: oData <= 16'h0000;
            14'h127a: oData <= 16'h0000;
            14'h127b: oData <= 16'h0000;
            14'h127c: oData <= 16'h8000;
            14'h127d: oData <= 16'h02aa;
            14'h127e: oData <= 16'h0000;
            14'h127f: oData <= 16'h0000;
            14'h1280: oData <= 16'h0000;
            14'h1281: oData <= 16'h0000;
            14'h1282: oData <= 16'h0a80;
            14'h1283: oData <= 16'h0000;
            14'h1284: oData <= 16'h0000;
            14'h1285: oData <= 16'h0000;
            14'h1286: oData <= 16'h0000;
            14'h1287: oData <= 16'h0000;
            14'h1288: oData <= 16'h0000;
            14'h1289: oData <= 16'h0000;
            14'h128a: oData <= 16'h0000;
            14'h128b: oData <= 16'h0000;
            14'h128c: oData <= 16'h0000;
            14'h128d: oData <= 16'h0000;
            14'h128e: oData <= 16'h0000;
            14'h128f: oData <= 16'h0000;
            14'h1290: oData <= 16'h0000;
            14'h1291: oData <= 16'h02aa;
            14'h1292: oData <= 16'h0000;
            14'h1293: oData <= 16'h0000;
            14'h1294: oData <= 16'h0000;
            14'h1295: oData <= 16'h0000;
            14'h1296: oData <= 16'h0000;
            14'h1297: oData <= 16'h0000;
            14'h1298: oData <= 16'h0000;
            14'h1299: oData <= 16'h0000;
            14'h129a: oData <= 16'h0000;
            14'h129b: oData <= 16'h0000;
            14'h129c: oData <= 16'h0000;
            14'h129d: oData <= 16'h0000;
            14'h129e: oData <= 16'h0000;
            14'h129f: oData <= 16'h0000;
            14'h12a0: oData <= 16'h0000;
            14'h12a1: oData <= 16'h0000;
            14'h12a2: oData <= 16'h0000;
            14'h12a3: oData <= 16'h0000;
            14'h12a4: oData <= 16'h0000;
            14'h12a5: oData <= 16'h02aa;
            14'h12a6: oData <= 16'h0000;
            14'h12a7: oData <= 16'h0000;
            14'h12a8: oData <= 16'h0000;
            14'h12a9: oData <= 16'h0000;
            14'h12aa: oData <= 16'h0000;
            14'h12ab: oData <= 16'h0000;
            14'h12ac: oData <= 16'h0000;
            14'h12ad: oData <= 16'h0000;
            14'h12ae: oData <= 16'h0000;
            14'h12af: oData <= 16'h0000;
            14'h12b0: oData <= 16'h0000;
            14'h12b1: oData <= 16'h0000;
            14'h12b2: oData <= 16'h0000;
            14'h12b3: oData <= 16'h0000;
            14'h12b4: oData <= 16'h0000;
            14'h12b5: oData <= 16'h0000;
            14'h12b6: oData <= 16'h0000;
            14'h12b7: oData <= 16'h0000;
            14'h12b8: oData <= 16'h0000;
            14'h12b9: oData <= 16'h00a8;
            14'h12ba: oData <= 16'h0000;
            14'h12bb: oData <= 16'h0000;
            14'h12bc: oData <= 16'h0000;
            14'h12bd: oData <= 16'h0000;
            14'h12be: oData <= 16'h0000;
            14'h12bf: oData <= 16'h0000;
            14'h12c0: oData <= 16'h0000;
            14'h12c1: oData <= 16'h0000;
            14'h12c2: oData <= 16'h0000;
            14'h12c3: oData <= 16'h0000;
            14'h12c4: oData <= 16'h0000;
            14'h12c5: oData <= 16'h0000;
            14'h12c6: oData <= 16'h0000;
            14'h12c7: oData <= 16'h0000;
            14'h12c8: oData <= 16'h0000;
            14'h12c9: oData <= 16'h0000;
            14'h12ca: oData <= 16'h0000;
            14'h12cb: oData <= 16'h0000;
            14'h12cc: oData <= 16'h0000;
            14'h12cd: oData <= 16'h0000;
            14'h12ce: oData <= 16'h0000;
            14'h12cf: oData <= 16'h0000;
            14'h12d0: oData <= 16'h0000;
            14'h12d1: oData <= 16'h0000;
            14'h12d2: oData <= 16'h0000;
            14'h12d3: oData <= 16'h000a;
            14'h12d4: oData <= 16'h0000;
            14'h12d5: oData <= 16'h0000;
            14'h12d6: oData <= 16'h0000;
            14'h12d7: oData <= 16'h0000;
            14'h12d8: oData <= 16'h0000;
            14'h12d9: oData <= 16'h0000;
            14'h12da: oData <= 16'h0000;
            14'h12db: oData <= 16'haaa8;
            14'h12dc: oData <= 16'haaaa;
            14'h12dd: oData <= 16'haaaa;
            14'h12de: oData <= 16'haaaa;
            14'h12df: oData <= 16'h02aa;
            14'h12e0: oData <= 16'h0000;
            14'h12e1: oData <= 16'h0000;
            14'h12e2: oData <= 16'h0000;
            14'h12e3: oData <= 16'h0000;
            14'h12e4: oData <= 16'h0000;
            14'h12e5: oData <= 16'h0000;
            14'h12e6: oData <= 16'h8000;
            14'h12e7: oData <= 16'h002a;
            14'h12e8: oData <= 16'h0000;
            14'h12e9: oData <= 16'h0000;
            14'h12ea: oData <= 16'h0000;
            14'h12eb: oData <= 16'h0000;
            14'h12ec: oData <= 16'h0000;
            14'h12ed: oData <= 16'h0000;
            14'h12ee: oData <= 16'h8000;
            14'h12ef: oData <= 16'haaaa;
            14'h12f0: oData <= 16'haaaa;
            14'h12f1: oData <= 16'haaaa;
            14'h12f2: oData <= 16'haaaa;
            14'h12f3: oData <= 16'haaaa;
            14'h12f4: oData <= 16'haaaa;
            14'h12f5: oData <= 16'h0000;
            14'h12f6: oData <= 16'h0000;
            14'h12f7: oData <= 16'h0000;
            14'h12f8: oData <= 16'h0000;
            14'h12f9: oData <= 16'h0000;
            14'h12fa: oData <= 16'h8000;
            14'h12fb: oData <= 16'h002a;
            14'h12fc: oData <= 16'h0000;
            14'h12fd: oData <= 16'h0000;
            14'h12fe: oData <= 16'h0000;
            14'h12ff: oData <= 16'h0000;
            14'h1300: oData <= 16'h0000;
            14'h1301: oData <= 16'h0000;
            14'h1302: oData <= 16'ha800;
            14'h1303: oData <= 16'hfffa;
            14'h1304: oData <= 16'hffff;
            14'h1305: oData <= 16'hffff;
            14'h1306: oData <= 16'hffff;
            14'h1307: oData <= 16'haaff;
            14'h1308: oData <= 16'haaaa;
            14'h1309: oData <= 16'h00aa;
            14'h130a: oData <= 16'h0000;
            14'h130b: oData <= 16'h0000;
            14'h130c: oData <= 16'h0000;
            14'h130d: oData <= 16'haa80;
            14'h130e: oData <= 16'h802a;
            14'h130f: oData <= 16'h002a;
            14'h1310: oData <= 16'h0000;
            14'h1311: oData <= 16'h0000;
            14'h1312: oData <= 16'h0000;
            14'h1313: oData <= 16'h0000;
            14'h1314: oData <= 16'h0000;
            14'h1315: oData <= 16'h0000;
            14'h1316: oData <= 16'haa00;
            14'h1317: oData <= 16'hffff;
            14'h1318: oData <= 16'hbfff;
            14'h1319: oData <= 16'haaaa;
            14'h131a: oData <= 16'haaaa;
            14'h131b: oData <= 16'hffff;
            14'h131c: oData <= 16'hbfff;
            14'h131d: oData <= 16'haaaa;
            14'h131e: oData <= 16'h0002;
            14'h131f: oData <= 16'h0000;
            14'h1320: oData <= 16'h0000;
            14'h1321: oData <= 16'haaa0;
            14'h1322: oData <= 16'h80aa;
            14'h1323: oData <= 16'h002a;
            14'h1324: oData <= 16'h0000;
            14'h1325: oData <= 16'h0000;
            14'h1326: oData <= 16'h0000;
            14'h1327: oData <= 16'h0000;
            14'h1328: oData <= 16'h0000;
            14'h1329: oData <= 16'h0000;
            14'h132a: oData <= 16'hfa80;
            14'h132b: oData <= 16'hffff;
            14'h132c: oData <= 16'heaff;
            14'h132d: oData <= 16'hffff;
            14'h132e: oData <= 16'hffff;
            14'h132f: oData <= 16'haaaa;
            14'h1330: oData <= 16'haaaa;
            14'h1331: oData <= 16'haabf;
            14'h1332: oData <= 16'h002a;
            14'h1333: oData <= 16'h0000;
            14'h1334: oData <= 16'h0000;
            14'h1335: oData <= 16'haaa8;
            14'h1336: oData <= 16'h82aa;
            14'h1337: oData <= 16'h002a;
            14'h1338: oData <= 16'h0000;
            14'h1339: oData <= 16'h0000;
            14'h133a: oData <= 16'h0000;
            14'h133b: oData <= 16'h0000;
            14'h133c: oData <= 16'h0000;
            14'h133d: oData <= 16'h0000;
            14'h133e: oData <= 16'hfea0;
            14'h133f: oData <= 16'hffff;
            14'h1340: oData <= 16'hffaf;
            14'h1341: oData <= 16'haaff;
            14'h1342: oData <= 16'hffea;
            14'h1343: oData <= 16'hffff;
            14'h1344: oData <= 16'hffff;
            14'h1345: oData <= 16'hffff;
            14'h1346: oData <= 16'h00aa;
            14'h1347: oData <= 16'h0000;
            14'h1348: oData <= 16'h0000;
            14'h1349: oData <= 16'haaa8;
            14'h134a: oData <= 16'h8aaa;
            14'h134b: oData <= 16'h002a;
            14'h134c: oData <= 16'h0000;
            14'h134d: oData <= 16'h0000;
            14'h134e: oData <= 16'h0000;
            14'h134f: oData <= 16'h0000;
            14'h1350: oData <= 16'h0000;
            14'h1351: oData <= 16'h0000;
            14'h1352: oData <= 16'hffa0;
            14'h1353: oData <= 16'hffff;
            14'h1354: oData <= 16'hbffa;
            14'h1355: oData <= 16'hffaa;
            14'h1356: oData <= 16'heabf;
            14'h1357: oData <= 16'hffff;
            14'h1358: oData <= 16'hffff;
            14'h1359: oData <= 16'hfaaa;
            14'h135a: oData <= 16'h0aaf;
            14'h135b: oData <= 16'h00a8;
            14'h135c: oData <= 16'h0000;
            14'h135d: oData <= 16'h02a8;
            14'h135e: oData <= 16'h8aa8;
            14'h135f: oData <= 16'h282a;
            14'h1360: oData <= 16'h0000;
            14'h1361: oData <= 16'h0000;
            14'h1362: oData <= 16'h0000;
            14'h1363: oData <= 16'h0000;
            14'h1364: oData <= 16'h0000;
            14'h1365: oData <= 16'h0000;
            14'h1366: oData <= 16'hffa8;
            14'h1367: oData <= 16'hafff;
            14'h1368: oData <= 16'heaff;
            14'h1369: oData <= 16'hffff;
            14'h136a: oData <= 16'hbfff;
            14'h136b: oData <= 16'haaaa;
            14'h136c: oData <= 16'haaaa;
            14'h136d: oData <= 16'hafff;
            14'h136e: oData <= 16'haabf;
            14'h136f: oData <= 16'h02aa;
            14'h1370: oData <= 16'h0000;
            14'h1371: oData <= 16'h02a8;
            14'h1372: oData <= 16'h8aa0;
            14'h1373: oData <= 16'haa2a;
            14'h1374: oData <= 16'h0000;
            14'h1375: oData <= 16'h0000;
            14'h1376: oData <= 16'h0000;
            14'h1377: oData <= 16'h0000;
            14'h1378: oData <= 16'h0000;
            14'h1379: oData <= 16'h0000;
            14'h137a: oData <= 16'hffea;
            14'h137b: oData <= 16'hfaff;
            14'h137c: oData <= 16'hffaf;
            14'h137d: oData <= 16'haaaf;
            14'h137e: oData <= 16'hffaa;
            14'h137f: oData <= 16'hffff;
            14'h1380: oData <= 16'hffff;
            14'h1381: oData <= 16'hbfff;
            14'h1382: oData <= 16'habff;
            14'h1383: oData <= 16'h02aa;
            14'h1384: oData <= 16'h0000;
            14'h1385: oData <= 16'h02a8;
            14'h1386: oData <= 16'h8aa0;
            14'h1387: oData <= 16'haaaa;
            14'h1388: oData <= 16'h0000;
            14'h1389: oData <= 16'h0000;
            14'h138a: oData <= 16'h0000;
            14'h138b: oData <= 16'h0000;
            14'h138c: oData <= 16'h0000;
            14'h138d: oData <= 16'h8000;
            14'h138e: oData <= 16'hfffa;
            14'h138f: oData <= 16'hffbf;
            14'h1390: oData <= 16'haffa;
            14'h1391: oData <= 16'hfffa;
            14'h1392: oData <= 16'hfebf;
            14'h1393: oData <= 16'hffff;
            14'h1394: oData <= 16'hbfff;
            14'h1395: oData <= 16'hffaa;
            14'h1396: oData <= 16'hbfff;
            14'h1397: oData <= 16'h00aa;
            14'h1398: oData <= 16'h0000;
            14'h1399: oData <= 16'h02a8;
            14'h139a: oData <= 16'h8aa0;
            14'h139b: oData <= 16'haaaa;
            14'h139c: oData <= 16'h0000;
            14'h139d: oData <= 16'h0000;
            14'h139e: oData <= 16'h0000;
            14'h139f: oData <= 16'h0000;
            14'h13a0: oData <= 16'h0000;
            14'h13a1: oData <= 16'h8000;
            14'h13a2: oData <= 16'hfffe;
            14'h13a3: oData <= 16'hafeb;
            14'h13a4: oData <= 16'hfabf;
            14'h13a5: oData <= 16'hffff;
            14'h13a6: oData <= 16'hffeb;
            14'h13a7: oData <= 16'hffff;
            14'h13a8: oData <= 16'heaaf;
            14'h13a9: oData <= 16'hfebf;
            14'h13aa: oData <= 16'hffff;
            14'h13ab: oData <= 16'h00aa;
            14'h13ac: oData <= 16'h0000;
            14'h13ad: oData <= 16'h02a8;
            14'h13ae: oData <= 16'h8aa0;
            14'h13af: oData <= 16'h2aaa;
            14'h13b0: oData <= 16'h0000;
            14'h13b1: oData <= 16'h0000;
            14'h13b2: oData <= 16'h0000;
            14'h13b3: oData <= 16'h0000;
            14'h13b4: oData <= 16'h0000;
            14'h13b5: oData <= 16'ha000;
            14'h13b6: oData <= 16'hfffe;
            14'h13b7: oData <= 16'hfbfe;
            14'h13b8: oData <= 16'hffeb;
            14'h13b9: oData <= 16'hffff;
            14'h13ba: oData <= 16'hffaf;
            14'h13bb: oData <= 16'hbfff;
            14'h13bc: oData <= 16'hfffa;
            14'h13bd: oData <= 16'hebff;
            14'h13be: oData <= 16'hffff;
            14'h13bf: oData <= 16'h02aa;
            14'h13c0: oData <= 16'h0000;
            14'h13c1: oData <= 16'h02a8;
            14'h13c2: oData <= 16'h8aa0;
            14'h13c3: oData <= 16'h02aa;
            14'h13c4: oData <= 16'h0000;
            14'h13c5: oData <= 16'h0000;
            14'h13c6: oData <= 16'h0000;
            14'h13c7: oData <= 16'h0000;
            14'h13c8: oData <= 16'h0000;
            14'h13c9: oData <= 16'ha000;
            14'h13ca: oData <= 16'hbfff;
            14'h13cb: oData <= 16'hfeff;
            14'h13cc: oData <= 16'hfffe;
            14'h13cd: oData <= 16'hffff;
            14'h13ce: oData <= 16'hffbf;
            14'h13cf: oData <= 16'hbfff;
            14'h13d0: oData <= 16'hffff;
            14'h13d1: oData <= 16'hbfff;
            14'h13d2: oData <= 16'hffff;
            14'h13d3: oData <= 16'h02aa;
            14'h13d4: oData <= 16'h0000;
            14'h13d5: oData <= 16'h2aa8;
            14'h13d6: oData <= 16'h0aa8;
            14'h13d7: oData <= 16'h00aa;
            14'h13d8: oData <= 16'h0000;
            14'h13d9: oData <= 16'h0000;
            14'h13da: oData <= 16'h0000;
            14'h13db: oData <= 16'h0000;
            14'h13dc: oData <= 16'h0000;
            14'h13dd: oData <= 16'ha000;
            14'h13de: oData <= 16'hffff;
            14'h13df: oData <= 16'hbfbf;
            14'h13e0: oData <= 16'hffff;
            14'h13e1: oData <= 16'hffff;
            14'h13e2: oData <= 16'hfebf;
            14'h13e3: oData <= 16'hffff;
            14'h13e4: oData <= 16'hffef;
            14'h13e5: oData <= 16'hbfff;
            14'h13e6: oData <= 16'hffff;
            14'h13e7: oData <= 16'h02ab;
            14'h13e8: oData <= 16'h0000;
            14'h13e9: oData <= 16'haaa8;
            14'h13ea: oData <= 16'h0aaa;
            14'h13eb: oData <= 16'h0000;
            14'h13ec: oData <= 16'h0000;
            14'h13ed: oData <= 16'h0000;
            14'h13ee: oData <= 16'h0000;
            14'h13ef: oData <= 16'h0000;
            14'h13f0: oData <= 16'h0000;
            14'h13f1: oData <= 16'ha800;
            14'h13f2: oData <= 16'hffff;
            14'h13f3: oData <= 16'hefef;
            14'h13f4: oData <= 16'hffff;
            14'h13f5: oData <= 16'hffff;
            14'h13f6: oData <= 16'hfeff;
            14'h13f7: oData <= 16'hffff;
            14'h13f8: oData <= 16'hfffb;
            14'h13f9: oData <= 16'hffff;
            14'h13fa: oData <= 16'hfffe;
            14'h13fb: oData <= 16'h02ab;
            14'h13fc: oData <= 16'h0000;
            14'h13fd: oData <= 16'haaa0;
            14'h13fe: oData <= 16'h02aa;
            14'h13ff: oData <= 16'h0000;
            14'h1400: oData <= 16'h0000;
            14'h1401: oData <= 16'h0000;
            14'h1402: oData <= 16'h0000;
            14'h1403: oData <= 16'h0000;
            14'h1404: oData <= 16'h0000;
            14'h1405: oData <= 16'he800;
            14'h1406: oData <= 16'hffff;
            14'h1407: oData <= 16'hfbff;
            14'h1408: oData <= 16'hafff;
            14'h1409: oData <= 16'hfeaa;
            14'h140a: oData <= 16'hfeff;
            14'h140b: oData <= 16'hffff;
            14'h140c: oData <= 16'hfffe;
            14'h140d: oData <= 16'hffff;
            14'h140e: oData <= 16'hfffe;
            14'h140f: oData <= 16'h0aab;
            14'h1410: oData <= 16'h0000;
            14'h1411: oData <= 16'haa80;
            14'h1412: oData <= 16'h02aa;
            14'h1413: oData <= 16'h0000;
            14'h1414: oData <= 16'h0000;
            14'h1415: oData <= 16'h0000;
            14'h1416: oData <= 16'h0000;
            14'h1417: oData <= 16'h0000;
            14'h1418: oData <= 16'h0000;
            14'h1419: oData <= 16'hea00;
            14'h141a: oData <= 16'hffff;
            14'h141b: oData <= 16'hffff;
            14'h141c: oData <= 16'haaaf;
            14'h141d: oData <= 16'haaaa;
            14'h141e: oData <= 16'hfeff;
            14'h141f: oData <= 16'hffff;
            14'h1420: oData <= 16'hfffe;
            14'h1421: oData <= 16'hffff;
            14'h1422: oData <= 16'hffff;
            14'h1423: oData <= 16'h0aab;
            14'h1424: oData <= 16'h0000;
            14'h1425: oData <= 16'ha800;
            14'h1426: oData <= 16'h002a;
            14'h1427: oData <= 16'h0000;
            14'h1428: oData <= 16'h0000;
            14'h1429: oData <= 16'h0000;
            14'h142a: oData <= 16'h0000;
            14'h142b: oData <= 16'h0000;
            14'h142c: oData <= 16'h0000;
            14'h142d: oData <= 16'hfa80;
            14'h142e: oData <= 16'hffff;
            14'h142f: oData <= 16'hffff;
            14'h1430: oData <= 16'haaaa;
            14'h1431: oData <= 16'haaea;
            14'h1432: oData <= 16'hfffa;
            14'h1433: oData <= 16'hffff;
            14'h1434: oData <= 16'hfffe;
            14'h1435: oData <= 16'hffff;
            14'h1436: oData <= 16'hffff;
            14'h1437: oData <= 16'h2aaf;
            14'h1438: oData <= 16'h0000;
            14'h1439: oData <= 16'h0000;
            14'h143a: oData <= 16'h0000;
            14'h143b: oData <= 16'h0000;
            14'h143c: oData <= 16'h0000;
            14'h143d: oData <= 16'h0000;
            14'h143e: oData <= 16'h0000;
            14'h143f: oData <= 16'h0000;
            14'h1440: oData <= 16'h0000;
            14'h1441: oData <= 16'hfea0;
            14'h1442: oData <= 16'hffff;
            14'h1443: oData <= 16'hbfff;
            14'h1444: oData <= 16'haaaa;
            14'h1445: oData <= 16'hbfea;
            14'h1446: oData <= 16'hffea;
            14'h1447: oData <= 16'hffff;
            14'h1448: oData <= 16'haafe;
            14'h1449: oData <= 16'hfaaa;
            14'h144a: oData <= 16'hffff;
            14'h144b: oData <= 16'h2aaf;
            14'h144c: oData <= 16'h0000;
            14'h144d: oData <= 16'h0000;
            14'h144e: oData <= 16'h0000;
            14'h144f: oData <= 16'h0000;
            14'h1450: oData <= 16'h0000;
            14'h1451: oData <= 16'h0000;
            14'h1452: oData <= 16'h0000;
            14'h1453: oData <= 16'h0000;
            14'h1454: oData <= 16'h0000;
            14'h1455: oData <= 16'haaa8;
            14'h1456: oData <= 16'hfffa;
            14'h1457: oData <= 16'hafaf;
            14'h1458: oData <= 16'haabe;
            14'h1459: oData <= 16'hffea;
            14'h145a: oData <= 16'hfeab;
            14'h145b: oData <= 16'hffff;
            14'h145c: oData <= 16'haaaf;
            14'h145d: oData <= 16'habff;
            14'h145e: oData <= 16'hffff;
            14'h145f: oData <= 16'haabf;
            14'h1460: oData <= 16'h0000;
            14'h1461: oData <= 16'h000a;
            14'h1462: oData <= 16'h0000;
            14'h1463: oData <= 16'h0000;
            14'h1464: oData <= 16'h0000;
            14'h1465: oData <= 16'h0000;
            14'h1466: oData <= 16'h0000;
            14'h1467: oData <= 16'h0000;
            14'h1468: oData <= 16'h0000;
            14'h1469: oData <= 16'hffaa;
            14'h146a: oData <= 16'hffff;
            14'h146b: oData <= 16'habfa;
            14'h146c: oData <= 16'haaaa;
            14'h146d: oData <= 16'hfeaa;
            14'h146e: oData <= 16'hfeaf;
            14'h146f: oData <= 16'hffff;
            14'h1470: oData <= 16'haaab;
            14'h1471: oData <= 16'haaaa;
            14'h1472: oData <= 16'hffef;
            14'h1473: oData <= 16'haabf;
            14'h1474: oData <= 16'ha800;
            14'h1475: oData <= 16'h002a;
            14'h1476: oData <= 16'h0000;
            14'h1477: oData <= 16'h0000;
            14'h1478: oData <= 16'h0000;
            14'h1479: oData <= 16'h0000;
            14'h147a: oData <= 16'h0000;
            14'h147b: oData <= 16'h0000;
            14'h147c: oData <= 16'h8000;
            14'h147d: oData <= 16'haaba;
            14'h147e: oData <= 16'hffaa;
            14'h147f: oData <= 16'habeb;
            14'h1480: oData <= 16'haaaa;
            14'h1481: oData <= 16'heaaa;
            14'h1482: oData <= 16'hfabf;
            14'h1483: oData <= 16'hebff;
            14'h1484: oData <= 16'haaaa;
            14'h1485: oData <= 16'haaaa;
            14'h1486: oData <= 16'habab;
            14'h1487: oData <= 16'haaea;
            14'h1488: oData <= 16'haa82;
            14'h1489: oData <= 16'h002a;
            14'h148a: oData <= 16'h0000;
            14'h148b: oData <= 16'h0000;
            14'h148c: oData <= 16'h0000;
            14'h148d: oData <= 16'h0000;
            14'h148e: oData <= 16'h0000;
            14'h148f: oData <= 16'h0000;
            14'h1490: oData <= 16'ha000;
            14'h1491: oData <= 16'hffee;
            14'h1492: oData <= 16'hffff;
            14'h1493: oData <= 16'hbebf;
            14'h1494: oData <= 16'hfffe;
            14'h1495: oData <= 16'haaff;
            14'h1496: oData <= 16'hfeaa;
            14'h1497: oData <= 16'haaff;
            14'h1498: oData <= 16'haaaa;
            14'h1499: oData <= 16'hfffe;
            14'h149a: oData <= 16'hfeff;
            14'h149b: oData <= 16'haabf;
            14'h149c: oData <= 16'haaaa;
            14'h149d: oData <= 16'h002a;
            14'h149e: oData <= 16'h0000;
            14'h149f: oData <= 16'h0000;
            14'h14a0: oData <= 16'h0000;
            14'h14a1: oData <= 16'h0000;
            14'h14a2: oData <= 16'h0000;
            14'h14a3: oData <= 16'h0000;
            14'h14a4: oData <= 16'ha800;
            14'h14a5: oData <= 16'hbffb;
            14'h14a6: oData <= 16'heaaa;
            14'h14a7: oData <= 16'hffbf;
            14'h14a8: oData <= 16'hafff;
            14'h14a9: oData <= 16'haffe;
            14'h14aa: oData <= 16'hfeaa;
            14'h14ab: oData <= 16'hafff;
            14'h14ac: oData <= 16'hffaa;
            14'h14ad: oData <= 16'hffff;
            14'h14ae: oData <= 16'hffff;
            14'h14af: oData <= 16'haafa;
            14'h14b0: oData <= 16'haaaa;
            14'h14b1: oData <= 16'h000a;
            14'h14b2: oData <= 16'h0000;
            14'h14b3: oData <= 16'h0000;
            14'h14b4: oData <= 16'h0000;
            14'h14b5: oData <= 16'h0000;
            14'h14b6: oData <= 16'h0000;
            14'h14b7: oData <= 16'h0000;
            14'h14b8: oData <= 16'hea00;
            14'h14b9: oData <= 16'habfe;
            14'h14ba: oData <= 16'haaaa;
            14'h14bb: oData <= 16'hfffa;
            14'h14bc: oData <= 16'habff;
            14'h14bd: oData <= 16'hffff;
            14'h14be: oData <= 16'hffeb;
            14'h14bf: oData <= 16'hffff;
            14'h14c0: oData <= 16'hfffa;
            14'h14c1: oData <= 16'hffff;
            14'h14c2: oData <= 16'hffff;
            14'h14c3: oData <= 16'habef;
            14'h14c4: oData <= 16'h2aaa;
            14'h14c5: oData <= 16'h0000;
            14'h14c6: oData <= 16'h0000;
            14'h14c7: oData <= 16'h0000;
            14'h14c8: oData <= 16'h0000;
            14'h14c9: oData <= 16'h0000;
            14'h14ca: oData <= 16'h0000;
            14'h14cb: oData <= 16'h0000;
            14'h14cc: oData <= 16'hba00;
            14'h14cd: oData <= 16'haaff;
            14'h14ce: oData <= 16'hafff;
            14'h14cf: oData <= 16'hffaa;
            14'h14d0: oData <= 16'heabf;
            14'h14d1: oData <= 16'hffff;
            14'h14d2: oData <= 16'hffff;
            14'h14d3: oData <= 16'hffff;
            14'h14d4: oData <= 16'hfffa;
            14'h14d5: oData <= 16'hffff;
            14'h14d6: oData <= 16'haaaf;
            14'h14d7: oData <= 16'hafbf;
            14'h14d8: oData <= 16'h02aa;
            14'h14d9: oData <= 16'h0000;
            14'h14da: oData <= 16'h0000;
            14'h14db: oData <= 16'h0000;
            14'h14dc: oData <= 16'h0000;
            14'h14dd: oData <= 16'h0000;
            14'h14de: oData <= 16'h0000;
            14'h14df: oData <= 16'h0000;
            14'h14e0: oData <= 16'hba80;
            14'h14e1: oData <= 16'hfaff;
            14'h14e2: oData <= 16'hfeff;
            14'h14e3: oData <= 16'haaaa;
            14'h14e4: oData <= 16'hfaaa;
            14'h14e5: oData <= 16'hffff;
            14'h14e6: oData <= 16'hffff;
            14'h14e7: oData <= 16'hffff;
            14'h14e8: oData <= 16'hfffa;
            14'h14e9: oData <= 16'hffff;
            14'h14ea: oData <= 16'haaab;
            14'h14eb: oData <= 16'hbfba;
            14'h14ec: oData <= 16'h000a;
            14'h14ed: oData <= 16'h0000;
            14'h14ee: oData <= 16'h0000;
            14'h14ef: oData <= 16'h0000;
            14'h14f0: oData <= 16'h0000;
            14'h14f1: oData <= 16'h0000;
            14'h14f2: oData <= 16'h0000;
            14'h14f3: oData <= 16'h0000;
            14'h14f4: oData <= 16'hbe80;
            14'h14f5: oData <= 16'hfabf;
            14'h14f6: oData <= 16'hfebf;
            14'h14f7: oData <= 16'haabf;
            14'h14f8: oData <= 16'hffaa;
            14'h14f9: oData <= 16'hffff;
            14'h14fa: oData <= 16'hffff;
            14'h14fb: oData <= 16'hffff;
            14'h14fc: oData <= 16'hfffa;
            14'h14fd: oData <= 16'hbfaf;
            14'h14fe: oData <= 16'hbfea;
            14'h14ff: oData <= 16'hbfba;
            14'h1500: oData <= 16'h000a;
            14'h1501: oData <= 16'h0000;
            14'h1502: oData <= 16'h0000;
            14'h1503: oData <= 16'h0000;
            14'h1504: oData <= 16'h0000;
            14'h1505: oData <= 16'h0000;
            14'h1506: oData <= 16'h0000;
            14'h1507: oData <= 16'h0000;
            14'h1508: oData <= 16'hbea0;
            14'h1509: oData <= 16'hfebf;
            14'h150a: oData <= 16'hfebf;
            14'h150b: oData <= 16'hffff;
            14'h150c: oData <= 16'hffff;
            14'h150d: oData <= 16'hffff;
            14'h150e: oData <= 16'hffff;
            14'h150f: oData <= 16'hffff;
            14'h1510: oData <= 16'hfffa;
            14'h1511: oData <= 16'haaaf;
            14'h1512: oData <= 16'hfffa;
            14'h1513: oData <= 16'hbfbb;
            14'h1514: oData <= 16'h000a;
            14'h1515: oData <= 16'h0000;
            14'h1516: oData <= 16'h0000;
            14'h1517: oData <= 16'h0000;
            14'h1518: oData <= 16'h0000;
            14'h1519: oData <= 16'h0000;
            14'h151a: oData <= 16'h0000;
            14'h151b: oData <= 16'h0000;
            14'h151c: oData <= 16'hbfa0;
            14'h151d: oData <= 16'hfeaf;
            14'h151e: oData <= 16'heabf;
            14'h151f: oData <= 16'hffff;
            14'h1520: oData <= 16'hffff;
            14'h1521: oData <= 16'hffff;
            14'h1522: oData <= 16'hffff;
            14'h1523: oData <= 16'hffff;
            14'h1524: oData <= 16'hffaa;
            14'h1525: oData <= 16'haabf;
            14'h1526: oData <= 16'hfefe;
            14'h1527: oData <= 16'hbeff;
            14'h1528: oData <= 16'h000a;
            14'h1529: oData <= 16'h0000;
            14'h152a: oData <= 16'h0000;
            14'h152b: oData <= 16'h0000;
            14'h152c: oData <= 16'h0000;
            14'h152d: oData <= 16'h0000;
            14'h152e: oData <= 16'h0000;
            14'h152f: oData <= 16'h0000;
            14'h1530: oData <= 16'hbfa0;
            14'h1531: oData <= 16'hffaf;
            14'h1532: oData <= 16'haaaf;
            14'h1533: oData <= 16'hfffe;
            14'h1534: oData <= 16'hffff;
            14'h1535: oData <= 16'hfbff;
            14'h1536: oData <= 16'hffaa;
            14'h1537: oData <= 16'hffff;
            14'h1538: oData <= 16'hfeab;
            14'h1539: oData <= 16'hffff;
            14'h153a: oData <= 16'hfebf;
            14'h153b: oData <= 16'hbeff;
            14'h153c: oData <= 16'h000a;
            14'h153d: oData <= 16'h0000;
            14'h153e: oData <= 16'h0000;
            14'h153f: oData <= 16'h0000;
            14'h1540: oData <= 16'h0000;
            14'h1541: oData <= 16'h0000;
            14'h1542: oData <= 16'h0000;
            14'h1543: oData <= 16'h0000;
            14'h1544: oData <= 16'hbfa0;
            14'h1545: oData <= 16'hffaf;
            14'h1546: oData <= 16'hafaa;
            14'h1547: oData <= 16'hffea;
            14'h1548: oData <= 16'hffff;
            14'h1549: oData <= 16'hbbff;
            14'h154a: oData <= 16'hfeaa;
            14'h154b: oData <= 16'hffff;
            14'h154c: oData <= 16'heabf;
            14'h154d: oData <= 16'hffff;
            14'h154e: oData <= 16'hfebf;
            14'h154f: oData <= 16'hbeff;
            14'h1550: oData <= 16'h000a;
            14'h1551: oData <= 16'h0000;
            14'h1552: oData <= 16'h0000;
            14'h1553: oData <= 16'h0000;
            14'h1554: oData <= 16'h0000;
            14'h1555: oData <= 16'h0000;
            14'h1556: oData <= 16'h0000;
            14'h1557: oData <= 16'h0000;
            14'h1558: oData <= 16'hbea0;
            14'h1559: oData <= 16'hafaf;
            14'h155a: oData <= 16'hffaa;
            14'h155b: oData <= 16'hfeaa;
            14'h155c: oData <= 16'habff;
            14'h155d: oData <= 16'haeaa;
            14'h155e: oData <= 16'hfffe;
            14'h155f: oData <= 16'hffff;
            14'h1560: oData <= 16'haaff;
            14'h1561: oData <= 16'hffff;
            14'h1562: oData <= 16'hfebf;
            14'h1563: oData <= 16'hefbf;
            14'h1564: oData <= 16'h000a;
            14'h1565: oData <= 16'h0000;
            14'h1566: oData <= 16'h0000;
            14'h1567: oData <= 16'h0000;
            14'h1568: oData <= 16'h0000;
            14'h1569: oData <= 16'h0000;
            14'h156a: oData <= 16'h0000;
            14'h156b: oData <= 16'h0000;
            14'h156c: oData <= 16'hbe80;
            14'h156d: oData <= 16'haeaf;
            14'h156e: oData <= 16'hfeae;
            14'h156f: oData <= 16'haaaf;
            14'h1570: oData <= 16'hfbff;
            14'h1571: oData <= 16'hafff;
            14'h1572: oData <= 16'hffff;
            14'h1573: oData <= 16'hffff;
            14'h1574: oData <= 16'haaff;
            14'h1575: oData <= 16'hfffe;
            14'h1576: oData <= 16'heabf;
            14'h1577: oData <= 16'hafeb;
            14'h1578: oData <= 16'h000a;
            14'h1579: oData <= 16'h0000;
            14'h157a: oData <= 16'h0000;
            14'h157b: oData <= 16'h0000;
            14'h157c: oData <= 16'h0000;
            14'h157d: oData <= 16'h0000;
            14'h157e: oData <= 16'h0000;
            14'h157f: oData <= 16'h0000;
            14'h1580: oData <= 16'hbe80;
            14'h1581: oData <= 16'hfebf;
            14'h1582: oData <= 16'hfebf;
            14'h1583: oData <= 16'haaff;
            14'h1584: oData <= 16'hfffa;
            14'h1585: oData <= 16'hafff;
            14'h1586: oData <= 16'haabf;
            14'h1587: oData <= 16'hfffa;
            14'h1588: oData <= 16'haabf;
            14'h1589: oData <= 16'hffeb;
            14'h158a: oData <= 16'heabf;
            14'h158b: oData <= 16'hbbff;
            14'h158c: oData <= 16'h0002;
            14'h158d: oData <= 16'h0000;
            14'h158e: oData <= 16'h0000;
            14'h158f: oData <= 16'h0000;
            14'h1590: oData <= 16'h0000;
            14'h1591: oData <= 16'h0000;
            14'h1592: oData <= 16'h0000;
            14'h1593: oData <= 16'h0000;
            14'h1594: oData <= 16'hfe80;
            14'h1595: oData <= 16'hfabe;
            14'h1596: oData <= 16'hfabf;
            14'h1597: oData <= 16'hafff;
            14'h1598: oData <= 16'hfeaa;
            14'h1599: oData <= 16'hafff;
            14'h159a: oData <= 16'haabe;
            14'h159b: oData <= 16'hfffa;
            14'h159c: oData <= 16'haebf;
            14'h159d: oData <= 16'hfebf;
            14'h159e: oData <= 16'heaaf;
            14'h159f: oData <= 16'hbeaf;
            14'h15a0: oData <= 16'h0002;
            14'h15a1: oData <= 16'h0000;
            14'h15a2: oData <= 16'h0000;
            14'h15a3: oData <= 16'h0000;
            14'h15a4: oData <= 16'h0000;
            14'h15a5: oData <= 16'h0000;
            14'h15a6: oData <= 16'h0000;
            14'h15a7: oData <= 16'h0000;
            14'h15a8: oData <= 16'hfa80;
            14'h15a9: oData <= 16'hfafe;
            14'h15aa: oData <= 16'heabf;
            14'h15ab: oData <= 16'hafff;
            14'h15ac: oData <= 16'haaab;
            14'h15ad: oData <= 16'hbffe;
            14'h15ae: oData <= 16'hffba;
            14'h15af: oData <= 16'hffff;
            14'h15b0: oData <= 16'hfeaf;
            14'h15b1: oData <= 16'hfbff;
            14'h15b2: oData <= 16'hebab;
            14'h15b3: oData <= 16'haffb;
            14'h15b4: oData <= 16'h0002;
            14'h15b5: oData <= 16'h0000;
            14'h15b6: oData <= 16'h0000;
            14'h15b7: oData <= 16'h0000;
            14'h15b8: oData <= 16'h0000;
            14'h15b9: oData <= 16'h0000;
            14'h15ba: oData <= 16'h0000;
            14'h15bb: oData <= 16'h0000;
            14'h15bc: oData <= 16'hea00;
            14'h15bd: oData <= 16'hfffb;
            14'h15be: oData <= 16'haabf;
            14'h15bf: oData <= 16'haffe;
            14'h15c0: oData <= 16'haaff;
            14'h15c1: oData <= 16'hffaa;
            14'h15c2: oData <= 16'hfffe;
            14'h15c3: oData <= 16'hebff;
            14'h15c4: oData <= 16'hffaa;
            14'h15c5: oData <= 16'hffff;
            14'h15c6: oData <= 16'heaaa;
            14'h15c7: oData <= 16'habff;
            14'h15c8: oData <= 16'h0000;
            14'h15c9: oData <= 16'h0000;
            14'h15ca: oData <= 16'h0000;
            14'h15cb: oData <= 16'h0000;
            14'h15cc: oData <= 16'h0000;
            14'h15cd: oData <= 16'h0000;
            14'h15ce: oData <= 16'h0000;
            14'h15cf: oData <= 16'h0000;
            14'h15d0: oData <= 16'he800;
            14'h15d1: oData <= 16'hffaf;
            14'h15d2: oData <= 16'haaff;
            14'h15d3: oData <= 16'hafea;
            14'h15d4: oData <= 16'hffff;
            14'h15d5: oData <= 16'heaaa;
            14'h15d6: oData <= 16'hffff;
            14'h15d7: oData <= 16'habff;
            14'h15d8: oData <= 16'hffea;
            14'h15d9: oData <= 16'hafff;
            14'h15da: oData <= 16'haaba;
            14'h15db: oData <= 16'h2bff;
            14'h15dc: oData <= 16'h0000;
            14'h15dd: oData <= 16'h0000;
            14'h15de: oData <= 16'h0000;
            14'h15df: oData <= 16'h0000;
            14'h15e0: oData <= 16'h0000;
            14'h15e1: oData <= 16'h0000;
            14'h15e2: oData <= 16'h0000;
            14'h15e3: oData <= 16'h0000;
            14'h15e4: oData <= 16'ha800;
            14'h15e5: oData <= 16'hfaff;
            14'h15e6: oData <= 16'habff;
            14'h15e7: oData <= 16'haeaa;
            14'h15e8: oData <= 16'hfffe;
            14'h15e9: oData <= 16'haabf;
            14'h15ea: oData <= 16'hffea;
            14'h15eb: oData <= 16'hafff;
            14'h15ec: oData <= 16'hfffe;
            14'h15ed: oData <= 16'haaff;
            14'h15ee: oData <= 16'haeba;
            14'h15ef: oData <= 16'h2aff;
            14'h15f0: oData <= 16'h0000;
            14'h15f1: oData <= 16'h0000;
            14'h15f2: oData <= 16'h0000;
            14'h15f3: oData <= 16'h0000;
            14'h15f4: oData <= 16'h0000;
            14'h15f5: oData <= 16'h0000;
            14'h15f6: oData <= 16'h0000;
            14'h15f7: oData <= 16'h0000;
            14'h15f8: oData <= 16'ha000;
            14'h15f9: oData <= 16'hffea;
            14'h15fa: oData <= 16'hafff;
            14'h15fb: oData <= 16'haaab;
            14'h15fc: oData <= 16'hfffa;
            14'h15fd: oData <= 16'haaff;
            14'h15fe: oData <= 16'haaaa;
            14'h15ff: oData <= 16'hfffe;
            14'h1600: oData <= 16'hffff;
            14'h1601: oData <= 16'heaab;
            14'h1602: oData <= 16'haaba;
            14'h1603: oData <= 16'h0aff;
            14'h1604: oData <= 16'h0000;
            14'h1605: oData <= 16'h0000;
            14'h1606: oData <= 16'h0000;
            14'h1607: oData <= 16'h0000;
            14'h1608: oData <= 16'h0000;
            14'h1609: oData <= 16'h0000;
            14'h160a: oData <= 16'h0000;
            14'h160b: oData <= 16'h0000;
            14'h160c: oData <= 16'h8000;
            14'h160d: oData <= 16'hffba;
            14'h160e: oData <= 16'hafff;
            14'h160f: oData <= 16'haafe;
            14'h1610: oData <= 16'hffea;
            14'h1611: oData <= 16'hfaff;
            14'h1612: oData <= 16'haaaf;
            14'h1613: oData <= 16'haaaa;
            14'h1614: oData <= 16'haaaa;
            14'h1615: oData <= 16'hfeaa;
            14'h1616: oData <= 16'haafa;
            14'h1617: oData <= 16'h0aff;
            14'h1618: oData <= 16'h0000;
            14'h1619: oData <= 16'h0000;
            14'h161a: oData <= 16'h0000;
            14'h161b: oData <= 16'h0000;
            14'h161c: oData <= 16'h0000;
            14'h161d: oData <= 16'h0000;
            14'h161e: oData <= 16'h0000;
            14'h161f: oData <= 16'h0000;
            14'h1620: oData <= 16'h0000;
            14'h1621: oData <= 16'hffea;
            14'h1622: oData <= 16'hbfff;
            14'h1623: oData <= 16'haffa;
            14'h1624: oData <= 16'hfaaa;
            14'h1625: oData <= 16'hfaff;
            14'h1626: oData <= 16'hffff;
            14'h1627: oData <= 16'haaaa;
            14'h1628: oData <= 16'haaaa;
            14'h1629: oData <= 16'hffaa;
            14'h162a: oData <= 16'haafa;
            14'h162b: oData <= 16'h0aff;
            14'h162c: oData <= 16'h0000;
            14'h162d: oData <= 16'h0000;
            14'h162e: oData <= 16'h0000;
            14'h162f: oData <= 16'h0000;
            14'h1630: oData <= 16'h0000;
            14'h1631: oData <= 16'h0000;
            14'h1632: oData <= 16'h0000;
            14'h1633: oData <= 16'h0000;
            14'h1634: oData <= 16'h0000;
            14'h1635: oData <= 16'hffa8;
            14'h1636: oData <= 16'hffff;
            14'h1637: oData <= 16'haffa;
            14'h1638: oData <= 16'haaaa;
            14'h1639: oData <= 16'hfabe;
            14'h163a: oData <= 16'hffff;
            14'h163b: oData <= 16'hfffa;
            14'h163c: oData <= 16'hffeb;
            14'h163d: oData <= 16'hfeaf;
            14'h163e: oData <= 16'haafa;
            14'h163f: oData <= 16'h0aff;
            14'h1640: oData <= 16'h0000;
            14'h1641: oData <= 16'h0000;
            14'h1642: oData <= 16'h0000;
            14'h1643: oData <= 16'h0000;
            14'h1644: oData <= 16'h0000;
            14'h1645: oData <= 16'h0000;
            14'h1646: oData <= 16'h0000;
            14'h1647: oData <= 16'h0000;
            14'h1648: oData <= 16'h0000;
            14'h1649: oData <= 16'hfea0;
            14'h164a: oData <= 16'hffff;
            14'h164b: oData <= 16'hafea;
            14'h164c: oData <= 16'haaaf;
            14'h164d: oData <= 16'hfeaa;
            14'h164e: oData <= 16'hffff;
            14'h164f: oData <= 16'hfffa;
            14'h1650: oData <= 16'hffeb;
            14'h1651: oData <= 16'hfebf;
            14'h1652: oData <= 16'haaba;
            14'h1653: oData <= 16'h0aff;
            14'h1654: oData <= 16'h0000;
            14'h1655: oData <= 16'h0000;
            14'h1656: oData <= 16'h0000;
            14'h1657: oData <= 16'h0000;
            14'h1658: oData <= 16'h0000;
            14'h1659: oData <= 16'h0000;
            14'h165a: oData <= 16'h0000;
            14'h165b: oData <= 16'h0000;
            14'h165c: oData <= 16'h0000;
            14'h165d: oData <= 16'hfa80;
            14'h165e: oData <= 16'hffff;
            14'h165f: oData <= 16'hafab;
            14'h1660: oData <= 16'haaff;
            14'h1661: oData <= 16'heaaa;
            14'h1662: oData <= 16'hffff;
            14'h1663: oData <= 16'hfffa;
            14'h1664: oData <= 16'hffeb;
            14'h1665: oData <= 16'hfebf;
            14'h1666: oData <= 16'haaaa;
            14'h1667: oData <= 16'h0aff;
            14'h1668: oData <= 16'h0000;
            14'h1669: oData <= 16'h0000;
            14'h166a: oData <= 16'h0000;
            14'h166b: oData <= 16'h0000;
            14'h166c: oData <= 16'h0000;
            14'h166d: oData <= 16'h0000;
            14'h166e: oData <= 16'h0000;
            14'h166f: oData <= 16'h0000;
            14'h1670: oData <= 16'h0000;
            14'h1671: oData <= 16'hfa00;
            14'h1672: oData <= 16'hffff;
            14'h1673: oData <= 16'haeaf;
            14'h1674: oData <= 16'hafff;
            14'h1675: oData <= 16'haaaa;
            14'h1676: oData <= 16'hffea;
            14'h1677: oData <= 16'hfffa;
            14'h1678: oData <= 16'hffeb;
            14'h1679: oData <= 16'haaaa;
            14'h167a: oData <= 16'haaaa;
            14'h167b: oData <= 16'h0aff;
            14'h167c: oData <= 16'h0000;
            14'h167d: oData <= 16'h0000;
            14'h167e: oData <= 16'h0000;
            14'h167f: oData <= 16'h0000;
            14'h1680: oData <= 16'h0000;
            14'h1681: oData <= 16'h0000;
            14'h1682: oData <= 16'h0000;
            14'h1683: oData <= 16'h0000;
            14'h1684: oData <= 16'h0000;
            14'h1685: oData <= 16'hfa00;
            14'h1686: oData <= 16'hffff;
            14'h1687: oData <= 16'haabf;
            14'h1688: oData <= 16'hffff;
            14'h1689: oData <= 16'haaaf;
            14'h168a: oData <= 16'haaaa;
            14'h168b: oData <= 16'haaaa;
            14'h168c: oData <= 16'haaaa;
            14'h168d: oData <= 16'haaaa;
            14'h168e: oData <= 16'haaaa;
            14'h168f: oData <= 16'h0aff;
            14'h1690: oData <= 16'h0000;
            14'h1691: oData <= 16'h0000;
            14'h1692: oData <= 16'h0000;
            14'h1693: oData <= 16'h0000;
            14'h1694: oData <= 16'h0000;
            14'h1695: oData <= 16'h0000;
            14'h1696: oData <= 16'h0000;
            14'h1697: oData <= 16'h0000;
            14'h1698: oData <= 16'h0000;
            14'h1699: oData <= 16'hea00;
            14'h169a: oData <= 16'hffff;
            14'h169b: oData <= 16'heaff;
            14'h169c: oData <= 16'hffff;
            14'h169d: oData <= 16'habaf;
            14'h169e: oData <= 16'haaaa;
            14'h169f: oData <= 16'haaaa;
            14'h16a0: oData <= 16'haaaa;
            14'h16a1: oData <= 16'haaaa;
            14'h16a2: oData <= 16'haaaa;
            14'h16a3: oData <= 16'h0aff;
            14'h16a4: oData <= 16'h0000;
            14'h16a5: oData <= 16'h0000;
            14'h16a6: oData <= 16'h0000;
            14'h16a7: oData <= 16'h0000;
            14'h16a8: oData <= 16'h0000;
            14'h16a9: oData <= 16'h0000;
            14'h16aa: oData <= 16'h0000;
            14'h16ab: oData <= 16'h0000;
            14'h16ac: oData <= 16'h0000;
            14'h16ad: oData <= 16'he800;
            14'h16ae: oData <= 16'hffff;
            14'h16af: oData <= 16'habff;
            14'h16b0: oData <= 16'hffff;
            14'h16b1: oData <= 16'hffaf;
            14'h16b2: oData <= 16'haaaa;
            14'h16b3: oData <= 16'haaaa;
            14'h16b4: oData <= 16'haaaa;
            14'h16b5: oData <= 16'haaaa;
            14'h16b6: oData <= 16'haaaa;
            14'h16b7: oData <= 16'h0aff;
            14'h16b8: oData <= 16'h0000;
            14'h16b9: oData <= 16'h0000;
            14'h16ba: oData <= 16'h0000;
            14'h16bb: oData <= 16'h0000;
            14'h16bc: oData <= 16'h0000;
            14'h16bd: oData <= 16'h0000;
            14'h16be: oData <= 16'h0000;
            14'h16bf: oData <= 16'h0000;
            14'h16c0: oData <= 16'h0000;
            14'h16c1: oData <= 16'ha800;
            14'h16c2: oData <= 16'hffff;
            14'h16c3: oData <= 16'hafff;
            14'h16c4: oData <= 16'hfffe;
            14'h16c5: oData <= 16'hffaf;
            14'h16c6: oData <= 16'haabf;
            14'h16c7: oData <= 16'haaaa;
            14'h16c8: oData <= 16'haaaa;
            14'h16c9: oData <= 16'haaaa;
            14'h16ca: oData <= 16'heaaa;
            14'h16cb: oData <= 16'h0aff;
            14'h16cc: oData <= 16'h0000;
            14'h16cd: oData <= 16'h0000;
            14'h16ce: oData <= 16'h0000;
            14'h16cf: oData <= 16'h0000;
            14'h16d0: oData <= 16'h0000;
            14'h16d1: oData <= 16'h0000;
            14'h16d2: oData <= 16'h0000;
            14'h16d3: oData <= 16'h0000;
            14'h16d4: oData <= 16'h0000;
            14'h16d5: oData <= 16'ha000;
            14'h16d6: oData <= 16'hfffe;
            14'h16d7: oData <= 16'hbfff;
            14'h16d8: oData <= 16'hffea;
            14'h16d9: oData <= 16'hffab;
            14'h16da: oData <= 16'hafff;
            14'h16db: oData <= 16'haaaa;
            14'h16dc: oData <= 16'haaaa;
            14'h16dd: oData <= 16'haaaa;
            14'h16de: oData <= 16'hebaa;
            14'h16df: oData <= 16'h0aff;
            14'h16e0: oData <= 16'h0000;
            14'h16e1: oData <= 16'h0000;
            14'h16e2: oData <= 16'h0000;
            14'h16e3: oData <= 16'h0000;
            14'h16e4: oData <= 16'h0000;
            14'h16e5: oData <= 16'h0000;
            14'h16e6: oData <= 16'h0000;
            14'h16e7: oData <= 16'h0000;
            14'h16e8: oData <= 16'h0000;
            14'h16e9: oData <= 16'h8000;
            14'h16ea: oData <= 16'hfffa;
            14'h16eb: oData <= 16'hffff;
            14'h16ec: oData <= 16'hffaa;
            14'h16ed: oData <= 16'hffeb;
            14'h16ee: oData <= 16'hafff;
            14'h16ef: oData <= 16'haabf;
            14'h16f0: oData <= 16'haaaa;
            14'h16f1: oData <= 16'haaaa;
            14'h16f2: oData <= 16'hebaf;
            14'h16f3: oData <= 16'h0aff;
            14'h16f4: oData <= 16'h0000;
            14'h16f5: oData <= 16'h0000;
            14'h16f6: oData <= 16'h0000;
            14'h16f7: oData <= 16'h0000;
            14'h16f8: oData <= 16'h0000;
            14'h16f9: oData <= 16'h0000;
            14'h16fa: oData <= 16'h0000;
            14'h16fb: oData <= 16'h0000;
            14'h16fc: oData <= 16'h0000;
            14'h16fd: oData <= 16'h0000;
            14'h16fe: oData <= 16'hffea;
            14'h16ff: oData <= 16'hffff;
            14'h1700: oData <= 16'hfaaf;
            14'h1701: oData <= 16'hffeb;
            14'h1702: oData <= 16'hafff;
            14'h1703: oData <= 16'hffff;
            14'h1704: oData <= 16'hffea;
            14'h1705: oData <= 16'hebfa;
            14'h1706: oData <= 16'hfaeb;
            14'h1707: oData <= 16'h0aff;
            14'h1708: oData <= 16'h0000;
            14'h1709: oData <= 16'h0000;
            14'h170a: oData <= 16'h0000;
            14'h170b: oData <= 16'h0000;
            14'h170c: oData <= 16'h0000;
            14'h170d: oData <= 16'h0000;
            14'h170e: oData <= 16'h0000;
            14'h170f: oData <= 16'h0000;
            14'h1710: oData <= 16'h0000;
            14'h1711: oData <= 16'h0000;
            14'h1712: oData <= 16'hffaa;
            14'h1713: oData <= 16'hffff;
            14'h1714: oData <= 16'haabf;
            14'h1715: oData <= 16'hffea;
            14'h1716: oData <= 16'hafff;
            14'h1717: oData <= 16'hffff;
            14'h1718: oData <= 16'hbffa;
            14'h1719: oData <= 16'heafa;
            14'h171a: oData <= 16'hfaaa;
            14'h171b: oData <= 16'h0aff;
            14'h171c: oData <= 16'h0000;
            14'h171d: oData <= 16'h0000;
            14'h171e: oData <= 16'h0000;
            14'h171f: oData <= 16'h0000;
            14'h1720: oData <= 16'h0000;
            14'h1721: oData <= 16'h0000;
            14'h1722: oData <= 16'h0000;
            14'h1723: oData <= 16'h0000;
            14'h1724: oData <= 16'h0000;
            14'h1725: oData <= 16'h0000;
            14'h1726: oData <= 16'hbea0;
            14'h1727: oData <= 16'hfaff;
            14'h1728: oData <= 16'habff;
            14'h1729: oData <= 16'hfffa;
            14'h172a: oData <= 16'hafff;
            14'h172b: oData <= 16'hffff;
            14'h172c: oData <= 16'hbffa;
            14'h172d: oData <= 16'hfafe;
            14'h172e: oData <= 16'hfebb;
            14'h172f: oData <= 16'h0aff;
            14'h1730: oData <= 16'h0000;
            14'h1731: oData <= 16'h0000;
            14'h1732: oData <= 16'h0000;
            14'h1733: oData <= 16'h0000;
            14'h1734: oData <= 16'h0000;
            14'h1735: oData <= 16'h0000;
            14'h1736: oData <= 16'h0000;
            14'h1737: oData <= 16'h0000;
            14'h1738: oData <= 16'h0000;
            14'h1739: oData <= 16'h0000;
            14'h173a: oData <= 16'hfa80;
            14'h173b: oData <= 16'hbffa;
            14'h173c: oData <= 16'hbfff;
            14'h173d: oData <= 16'hfeaa;
            14'h173e: oData <= 16'hafff;
            14'h173f: oData <= 16'hffff;
            14'h1740: oData <= 16'haffa;
            14'h1741: oData <= 16'hfabe;
            14'h1742: oData <= 16'hfeaf;
            14'h1743: oData <= 16'h0aff;
            14'h1744: oData <= 16'h0000;
            14'h1745: oData <= 16'h0000;
            14'h1746: oData <= 16'h0000;
            14'h1747: oData <= 16'h0000;
            14'h1748: oData <= 16'h0000;
            14'h1749: oData <= 16'h0000;
            14'h174a: oData <= 16'h0000;
            14'h174b: oData <= 16'h0000;
            14'h174c: oData <= 16'h0000;
            14'h174d: oData <= 16'h0000;
            14'h174e: oData <= 16'hea00;
            14'h174f: oData <= 16'hffaf;
            14'h1750: oData <= 16'hfffa;
            14'h1751: oData <= 16'haaab;
            14'h1752: oData <= 16'hafff;
            14'h1753: oData <= 16'hbfff;
            14'h1754: oData <= 16'haffa;
            14'h1755: oData <= 16'haaff;
            14'h1756: oData <= 16'hffea;
            14'h1757: oData <= 16'h0aff;
            14'h1758: oData <= 16'h0000;
            14'h1759: oData <= 16'h0000;
            14'h175a: oData <= 16'h0000;
            14'h175b: oData <= 16'h0000;
            14'h175c: oData <= 16'h0000;
            14'h175d: oData <= 16'h0000;
            14'h175e: oData <= 16'h0000;
            14'h175f: oData <= 16'h0000;
            14'h1760: oData <= 16'h0000;
            14'h1761: oData <= 16'h0000;
            14'h1762: oData <= 16'ha800;
            14'h1763: oData <= 16'hfafe;
            14'h1764: oData <= 16'hffaf;
            14'h1765: oData <= 16'haaff;
            14'h1766: oData <= 16'haaaa;
            14'h1767: oData <= 16'hbffe;
            14'h1768: oData <= 16'habfe;
            14'h1769: oData <= 16'haaaa;
            14'h176a: oData <= 16'hfffa;
            14'h176b: oData <= 16'h0aff;
            14'h176c: oData <= 16'h0000;
            14'h176d: oData <= 16'h0000;
            14'h176e: oData <= 16'h0000;
            14'h176f: oData <= 16'h0000;
            14'h1770: oData <= 16'h0000;
            14'h1771: oData <= 16'h0000;
            14'h1772: oData <= 16'h0000;
            14'h1773: oData <= 16'h0000;
            14'h1774: oData <= 16'h0000;
            14'h1775: oData <= 16'h0000;
            14'h1776: oData <= 16'ha000;
            14'h1777: oData <= 16'haffa;
            14'h1778: oData <= 16'hfaff;
            14'h1779: oData <= 16'hbfff;
            14'h177a: oData <= 16'haaaa;
            14'h177b: oData <= 16'haaaa;
            14'h177c: oData <= 16'haaaa;
            14'h177d: oData <= 16'hfaaa;
            14'h177e: oData <= 16'hffff;
            14'h177f: oData <= 16'h0aff;
            14'h1780: oData <= 16'h0000;
            14'h1781: oData <= 16'h0000;
            14'h1782: oData <= 16'h0000;
            14'h1783: oData <= 16'h0000;
            14'h1784: oData <= 16'h0000;
            14'h1785: oData <= 16'h0000;
            14'h1786: oData <= 16'h0000;
            14'h1787: oData <= 16'h0000;
            14'h1788: oData <= 16'h0000;
            14'h1789: oData <= 16'h0000;
            14'h178a: oData <= 16'h0000;
            14'h178b: oData <= 16'hffaa;
            14'h178c: oData <= 16'haffa;
            14'h178d: oData <= 16'hffff;
            14'h178e: oData <= 16'hffff;
            14'h178f: oData <= 16'haaaa;
            14'h1790: oData <= 16'hfaaa;
            14'h1791: oData <= 16'hffff;
            14'h1792: oData <= 16'hffff;
            14'h1793: oData <= 16'h0aff;
            14'h1794: oData <= 16'h0000;
            14'h1795: oData <= 16'h0000;
            14'h1796: oData <= 16'h0000;
            14'h1797: oData <= 16'h0000;
            14'h1798: oData <= 16'h0000;
            14'h1799: oData <= 16'h0000;
            14'h179a: oData <= 16'h0000;
            14'h179b: oData <= 16'h0000;
            14'h179c: oData <= 16'h0000;
            14'h179d: oData <= 16'h0000;
            14'h179e: oData <= 16'h0000;
            14'h179f: oData <= 16'hfaa8;
            14'h17a0: oData <= 16'hffaf;
            14'h17a1: oData <= 16'hffea;
            14'h17a2: oData <= 16'hffff;
            14'h17a3: oData <= 16'hffff;
            14'h17a4: oData <= 16'hffff;
            14'h17a5: oData <= 16'hffff;
            14'h17a6: oData <= 16'hffbf;
            14'h17a7: oData <= 16'h2aff;
            14'h17a8: oData <= 16'h0000;
            14'h17a9: oData <= 16'h0000;
            14'h17aa: oData <= 16'h0000;
            14'h17ab: oData <= 16'h0000;
            14'h17ac: oData <= 16'h0000;
            14'h17ad: oData <= 16'h0000;
            14'h17ae: oData <= 16'h0000;
            14'h17af: oData <= 16'h0000;
            14'h17b0: oData <= 16'h0000;
            14'h17b1: oData <= 16'h0000;
            14'h17b2: oData <= 16'h0000;
            14'h17b3: oData <= 16'haa80;
            14'h17b4: oData <= 16'hfaff;
            14'h17b5: oData <= 16'hfabf;
            14'h17b6: oData <= 16'hffff;
            14'h17b7: oData <= 16'hffff;
            14'h17b8: oData <= 16'hffff;
            14'h17b9: oData <= 16'hffff;
            14'h17ba: oData <= 16'hbfef;
            14'h17bb: oData <= 16'h2bff;
            14'h17bc: oData <= 16'h0000;
            14'h17bd: oData <= 16'h0000;
            14'h17be: oData <= 16'h0000;
            14'h17bf: oData <= 16'h0000;
            14'h17c0: oData <= 16'h0000;
            14'h17c1: oData <= 16'h0000;
            14'h17c2: oData <= 16'h0000;
            14'h17c3: oData <= 16'h0000;
            14'h17c4: oData <= 16'h0000;
            14'h17c5: oData <= 16'h0000;
            14'h17c6: oData <= 16'h0000;
            14'h17c7: oData <= 16'ha800;
            14'h17c8: oData <= 16'haffa;
            14'h17c9: oData <= 16'haffe;
            14'h17ca: oData <= 16'hffff;
            14'h17cb: oData <= 16'haaaa;
            14'h17cc: oData <= 16'haaaa;
            14'h17cd: oData <= 16'hffff;
            14'h17ce: oData <= 16'hbffa;
            14'h17cf: oData <= 16'h2bff;
            14'h17d0: oData <= 16'h0000;
            14'h17d1: oData <= 16'h0000;
            14'h17d2: oData <= 16'h0000;
            14'h17d3: oData <= 16'h0000;
            14'h17d4: oData <= 16'h0000;
            14'h17d5: oData <= 16'h0000;
            14'h17d6: oData <= 16'h0000;
            14'h17d7: oData <= 16'h0000;
            14'h17d8: oData <= 16'h0000;
            14'h17d9: oData <= 16'h0000;
            14'h17da: oData <= 16'h0000;
            14'h17db: oData <= 16'h8000;
            14'h17dc: oData <= 16'hffaa;
            14'h17dd: oData <= 16'hffab;
            14'h17de: oData <= 16'hfeaa;
            14'h17df: oData <= 16'hffff;
            14'h17e0: oData <= 16'hffff;
            14'h17e1: oData <= 16'hbfff;
            14'h17e2: oData <= 16'hbfff;
            14'h17e3: oData <= 16'h2bff;
            14'h17e4: oData <= 16'h0000;
            14'h17e5: oData <= 16'h0000;
            14'h17e6: oData <= 16'h0000;
            14'h17e7: oData <= 16'h0000;
            14'h17e8: oData <= 16'h0000;
            14'h17e9: oData <= 16'h0a00;
            14'h17ea: oData <= 16'h0000;
            14'h17eb: oData <= 16'h0000;
            14'h17ec: oData <= 16'h0000;
            14'h17ed: oData <= 16'h0000;
            14'h17ee: oData <= 16'h0000;
            14'h17ef: oData <= 16'h0000;
            14'h17f0: oData <= 16'heaa8;
            14'h17f1: oData <= 16'heaff;
            14'h17f2: oData <= 16'habff;
            14'h17f3: oData <= 16'haaaa;
            14'h17f4: oData <= 16'hffff;
            14'h17f5: oData <= 16'heabf;
            14'h17f6: oData <= 16'hefff;
            14'h17f7: oData <= 16'h2bff;
            14'h17f8: oData <= 16'h0000;
            14'h17f9: oData <= 16'h0000;
            14'h17fa: oData <= 16'h0000;
            14'h17fb: oData <= 16'h0000;
            14'h17fc: oData <= 16'h0000;
            14'h17fd: oData <= 16'h2a80;
            14'h17fe: oData <= 16'h0000;
            14'h17ff: oData <= 16'h0000;
            14'h1800: oData <= 16'h0000;
            14'h1801: oData <= 16'h0000;
            14'h1802: oData <= 16'h0000;
            14'h1803: oData <= 16'h0000;
            14'h1804: oData <= 16'haa80;
            14'h1805: oData <= 16'hbffe;
            14'h1806: oData <= 16'hffaa;
            14'h1807: oData <= 16'hffff;
            14'h1808: oData <= 16'haaaa;
            14'h1809: oData <= 16'hffea;
            14'h180a: oData <= 16'hfaff;
            14'h180b: oData <= 16'h2bff;
            14'h180c: oData <= 16'h0000;
            14'h180d: oData <= 16'h0000;
            14'h180e: oData <= 16'h0000;
            14'h180f: oData <= 16'h0000;
            14'h1810: oData <= 16'h0000;
            14'h1811: oData <= 16'h2aa0;
            14'h1812: oData <= 16'h0000;
            14'h1813: oData <= 16'h0000;
            14'h1814: oData <= 16'h0000;
            14'h1815: oData <= 16'h0000;
            14'h1816: oData <= 16'h0000;
            14'h1817: oData <= 16'h0000;
            14'h1818: oData <= 16'ha000;
            14'h1819: oData <= 16'hffea;
            14'h181a: oData <= 16'haaff;
            14'h181b: oData <= 16'hfffa;
            14'h181c: oData <= 16'hffff;
            14'h181d: oData <= 16'hffff;
            14'h181e: oData <= 16'hffbf;
            14'h181f: oData <= 16'h2bff;
            14'h1820: oData <= 16'h0000;
            14'h1821: oData <= 16'h0000;
            14'h1822: oData <= 16'h0000;
            14'h1823: oData <= 16'h0000;
            14'h1824: oData <= 16'h0000;
            14'h1825: oData <= 16'h2aa0;
            14'h1826: oData <= 16'h0000;
            14'h1827: oData <= 16'h0000;
            14'h1828: oData <= 16'h0000;
            14'h1829: oData <= 16'h0000;
            14'h182a: oData <= 16'h0000;
            14'h182b: oData <= 16'h0000;
            14'h182c: oData <= 16'h0000;
            14'h182d: oData <= 16'hfeaa;
            14'h182e: oData <= 16'hffff;
            14'h182f: oData <= 16'haaaf;
            14'h1830: oData <= 16'hffaa;
            14'h1831: oData <= 16'hbfff;
            14'h1832: oData <= 16'hffea;
            14'h1833: oData <= 16'h2aff;
            14'h1834: oData <= 16'h0000;
            14'h1835: oData <= 16'h0000;
            14'h1836: oData <= 16'h0000;
            14'h1837: oData <= 16'h0000;
            14'h1838: oData <= 16'h0000;
            14'h1839: oData <= 16'h0aa8;
            14'h183a: oData <= 16'h0000;
            14'h183b: oData <= 16'h0000;
            14'h183c: oData <= 16'h0000;
            14'h183d: oData <= 16'h0000;
            14'h183e: oData <= 16'h0000;
            14'h183f: oData <= 16'h0000;
            14'h1840: oData <= 16'h0000;
            14'h1841: oData <= 16'heaa0;
            14'h1842: oData <= 16'hffff;
            14'h1843: oData <= 16'hffff;
            14'h1844: oData <= 16'haaff;
            14'h1845: oData <= 16'heaaa;
            14'h1846: oData <= 16'hffff;
            14'h1847: oData <= 16'h0aff;
            14'h1848: oData <= 16'h0000;
            14'h1849: oData <= 16'h0000;
            14'h184a: oData <= 16'h0000;
            14'h184b: oData <= 16'h0000;
            14'h184c: oData <= 16'h0000;
            14'h184d: oData <= 16'h0aa8;
            14'h184e: oData <= 16'h0000;
            14'h184f: oData <= 16'h0000;
            14'h1850: oData <= 16'h0000;
            14'h1851: oData <= 16'h0000;
            14'h1852: oData <= 16'h0000;
            14'h1853: oData <= 16'h0000;
            14'h1854: oData <= 16'h0000;
            14'h1855: oData <= 16'haa00;
            14'h1856: oData <= 16'hfffe;
            14'h1857: oData <= 16'hffff;
            14'h1858: oData <= 16'hffff;
            14'h1859: oData <= 16'hffff;
            14'h185a: oData <= 16'hffff;
            14'h185b: oData <= 16'h0abf;
            14'h185c: oData <= 16'h0000;
            14'h185d: oData <= 16'h0000;
            14'h185e: oData <= 16'h0000;
            14'h185f: oData <= 16'h0000;
            14'h1860: oData <= 16'h0000;
            14'h1861: oData <= 16'h02aa;
            14'h1862: oData <= 16'h0000;
            14'h1863: oData <= 16'h0000;
            14'h1864: oData <= 16'h0000;
            14'h1865: oData <= 16'h0000;
            14'h1866: oData <= 16'h0000;
            14'h1867: oData <= 16'h0000;
            14'h1868: oData <= 16'h0000;
            14'h1869: oData <= 16'ha000;
            14'h186a: oData <= 16'hffea;
            14'h186b: oData <= 16'hffff;
            14'h186c: oData <= 16'hffff;
            14'h186d: oData <= 16'hffff;
            14'h186e: oData <= 16'hffff;
            14'h186f: oData <= 16'h02bf;
            14'h1870: oData <= 16'h0000;
            14'h1871: oData <= 16'h0000;
            14'h1872: oData <= 16'h0000;
            14'h1873: oData <= 16'h0000;
            14'h1874: oData <= 16'h0000;
            14'h1875: oData <= 16'h02aa;
            14'h1876: oData <= 16'h0000;
            14'h1877: oData <= 16'h0000;
            14'h1878: oData <= 16'h0000;
            14'h1879: oData <= 16'h0000;
            14'h187a: oData <= 16'h0000;
            14'h187b: oData <= 16'h0000;
            14'h187c: oData <= 16'h0000;
            14'h187d: oData <= 16'h0000;
            14'h187e: oData <= 16'haaaa;
            14'h187f: oData <= 16'hffff;
            14'h1880: oData <= 16'hffff;
            14'h1881: oData <= 16'hffff;
            14'h1882: oData <= 16'hffff;
            14'h1883: oData <= 16'h02af;
            14'h1884: oData <= 16'h0000;
            14'h1885: oData <= 16'h0000;
            14'h1886: oData <= 16'h0000;
            14'h1887: oData <= 16'h0000;
            14'h1888: oData <= 16'h0000;
            14'h1889: oData <= 16'h00aa;
            14'h188a: oData <= 16'h0000;
            14'h188b: oData <= 16'h02a8;
            14'h188c: oData <= 16'h0000;
            14'h188d: oData <= 16'h0000;
            14'h188e: oData <= 16'h0000;
            14'h188f: oData <= 16'h0000;
            14'h1890: oData <= 16'h0000;
            14'h1891: oData <= 16'h0000;
            14'h1892: oData <= 16'haaa0;
            14'h1893: oData <= 16'hffaa;
            14'h1894: oData <= 16'hffff;
            14'h1895: oData <= 16'hffff;
            14'h1896: oData <= 16'hffff;
            14'h1897: oData <= 16'h00aa;
            14'h1898: oData <= 16'h0000;
            14'h1899: oData <= 16'h0000;
            14'h189a: oData <= 16'h0000;
            14'h189b: oData <= 16'h0000;
            14'h189c: oData <= 16'h8000;
            14'h189d: oData <= 16'h00aa;
            14'h189e: oData <= 16'h0000;
            14'h189f: oData <= 16'h0aaa;
            14'h18a0: oData <= 16'h0000;
            14'h18a1: oData <= 16'h0000;
            14'h18a2: oData <= 16'h0000;
            14'h18a3: oData <= 16'h0000;
            14'h18a4: oData <= 16'h0000;
            14'h18a5: oData <= 16'h0000;
            14'h18a6: oData <= 16'haa80;
            14'h18a7: oData <= 16'haaaa;
            14'h18a8: oData <= 16'hffff;
            14'h18a9: oData <= 16'hffff;
            14'h18aa: oData <= 16'hbfff;
            14'h18ab: oData <= 16'h002a;
            14'h18ac: oData <= 16'h0000;
            14'h18ad: oData <= 16'h0000;
            14'h18ae: oData <= 16'h0000;
            14'h18af: oData <= 16'h0000;
            14'h18b0: oData <= 16'h8000;
            14'h18b1: oData <= 16'h00aa;
            14'h18b2: oData <= 16'h8000;
            14'h18b3: oData <= 16'h0aaa;
            14'h18b4: oData <= 16'h0000;
            14'h18b5: oData <= 16'h0000;
            14'h18b6: oData <= 16'h0000;
            14'h18b7: oData <= 16'h0000;
            14'h18b8: oData <= 16'h0000;
            14'h18b9: oData <= 16'h0000;
            14'h18ba: oData <= 16'haa80;
            14'h18bb: oData <= 16'haa82;
            14'h18bc: oData <= 16'hffaa;
            14'h18bd: oData <= 16'hffff;
            14'h18be: oData <= 16'haaff;
            14'h18bf: oData <= 16'h0002;
            14'h18c0: oData <= 16'h0000;
            14'h18c1: oData <= 16'h0000;
            14'h18c2: oData <= 16'h0000;
            14'h18c3: oData <= 16'h0000;
            14'h18c4: oData <= 16'h8000;
            14'h18c5: oData <= 16'h002a;
            14'h18c6: oData <= 16'ha000;
            14'h18c7: oData <= 16'h2aaa;
            14'h18c8: oData <= 16'h0000;
            14'h18c9: oData <= 16'h0000;
            14'h18ca: oData <= 16'h0000;
            14'h18cb: oData <= 16'h0000;
            14'h18cc: oData <= 16'h0000;
            14'h18cd: oData <= 16'h0000;
            14'h18ce: oData <= 16'haa00;
            14'h18cf: oData <= 16'ha002;
            14'h18d0: oData <= 16'haaaa;
            14'h18d1: oData <= 16'haaaa;
            14'h18d2: oData <= 16'h2aaa;
            14'h18d3: oData <= 16'h0000;
            14'h18d4: oData <= 16'h0000;
            14'h18d5: oData <= 16'h0000;
            14'h18d6: oData <= 16'h0000;
            14'h18d7: oData <= 16'h0000;
            14'h18d8: oData <= 16'ha000;
            14'h18d9: oData <= 16'h002a;
            14'h18da: oData <= 16'ha800;
            14'h18db: oData <= 16'h2aaa;
            14'h18dc: oData <= 16'h0000;
            14'h18dd: oData <= 16'h0000;
            14'h18de: oData <= 16'h0000;
            14'h18df: oData <= 16'h0000;
            14'h18e0: oData <= 16'h0000;
            14'h18e1: oData <= 16'h0000;
            14'h18e2: oData <= 16'haa00;
            14'h18e3: oData <= 16'ha802;
            14'h18e4: oData <= 16'haaaa;
            14'h18e5: oData <= 16'haaaa;
            14'h18e6: oData <= 16'h02aa;
            14'h18e7: oData <= 16'h0000;
            14'h18e8: oData <= 16'h0000;
            14'h18e9: oData <= 16'h0000;
            14'h18ea: oData <= 16'h0000;
            14'h18eb: oData <= 16'h0000;
            14'h18ec: oData <= 16'ha000;
            14'h18ed: oData <= 16'h002a;
            14'h18ee: oData <= 16'ha800;
            14'h18ef: oData <= 16'h2a8a;
            14'h18f0: oData <= 16'h2800;
            14'h18f1: oData <= 16'h0000;
            14'h18f2: oData <= 16'h0000;
            14'h18f3: oData <= 16'h0000;
            14'h18f4: oData <= 16'h0000;
            14'h18f5: oData <= 16'h0000;
            14'h18f6: oData <= 16'haa00;
            14'h18f7: oData <= 16'ha802;
            14'h18f8: oData <= 16'h000a;
            14'h18f9: oData <= 16'haaaa;
            14'h18fa: oData <= 16'h0aaa;
            14'h18fb: oData <= 16'h0000;
            14'h18fc: oData <= 16'h0000;
            14'h18fd: oData <= 16'h0000;
            14'h18fe: oData <= 16'h0000;
            14'h18ff: oData <= 16'h0000;
            14'h1900: oData <= 16'ha000;
            14'h1901: oData <= 16'h000a;
            14'h1902: oData <= 16'ha800;
            14'h1903: oData <= 16'h2a82;
            14'h1904: oData <= 16'haa00;
            14'h1905: oData <= 16'h0000;
            14'h1906: oData <= 16'h0000;
            14'h1907: oData <= 16'h0000;
            14'h1908: oData <= 16'h0000;
            14'h1909: oData <= 16'h0000;
            14'h190a: oData <= 16'haa00;
            14'h190b: oData <= 16'haa0a;
            14'h190c: oData <= 16'h000a;
            14'h190d: oData <= 16'haa80;
            14'h190e: oData <= 16'h0aaa;
            14'h190f: oData <= 16'h0000;
            14'h1910: oData <= 16'h0000;
            14'h1911: oData <= 16'h0000;
            14'h1912: oData <= 16'h0000;
            14'h1913: oData <= 16'h0000;
            14'h1914: oData <= 16'ha000;
            14'h1915: oData <= 16'h000a;
            14'h1916: oData <= 16'haa00;
            14'h1917: oData <= 16'h2a82;
            14'h1918: oData <= 16'haa80;
            14'h1919: oData <= 16'h0000;
            14'h191a: oData <= 16'h0000;
            14'h191b: oData <= 16'h0000;
            14'h191c: oData <= 16'h0000;
            14'h191d: oData <= 16'h0000;
            14'h191e: oData <= 16'ha800;
            14'h191f: oData <= 16'haa8a;
            14'h1920: oData <= 16'h0002;
            14'h1921: oData <= 16'ha800;
            14'h1922: oData <= 16'h0aaa;
            14'h1923: oData <= 16'h0000;
            14'h1924: oData <= 16'h0000;
            14'h1925: oData <= 16'h0000;
            14'h1926: oData <= 16'h0000;
            14'h1927: oData <= 16'h0000;
            14'h1928: oData <= 16'ha000;
            14'h1929: oData <= 16'h002a;
            14'h192a: oData <= 16'haa00;
            14'h192b: oData <= 16'h2a82;
            14'h192c: oData <= 16'haa80;
            14'h192d: oData <= 16'h0000;
            14'h192e: oData <= 16'h0000;
            14'h192f: oData <= 16'h0000;
            14'h1930: oData <= 16'h0000;
            14'h1931: oData <= 16'h0000;
            14'h1932: oData <= 16'ha800;
            14'h1933: oData <= 16'haaaa;
            14'h1934: oData <= 16'h0000;
            14'h1935: oData <= 16'h0000;
            14'h1936: oData <= 16'h02aa;
            14'h1937: oData <= 16'h0000;
            14'h1938: oData <= 16'h0000;
            14'h1939: oData <= 16'h0000;
            14'h193a: oData <= 16'h0000;
            14'h193b: oData <= 16'h0000;
            14'h193c: oData <= 16'ha000;
            14'h193d: oData <= 16'h00aa;
            14'h193e: oData <= 16'haa00;
            14'h193f: oData <= 16'h2a80;
            14'h1940: oData <= 16'h2aa0;
            14'h1941: oData <= 16'h0000;
            14'h1942: oData <= 16'h0000;
            14'h1943: oData <= 16'h0000;
            14'h1944: oData <= 16'h0000;
            14'h1945: oData <= 16'h0000;
            14'h1946: oData <= 16'ha800;
            14'h1947: oData <= 16'h2aaa;
            14'h1948: oData <= 16'h0000;
            14'h1949: oData <= 16'h0000;
            14'h194a: oData <= 16'h0000;
            14'h194b: oData <= 16'h0000;
            14'h194c: oData <= 16'h0000;
            14'h194d: oData <= 16'h0000;
            14'h194e: oData <= 16'h0000;
            14'h194f: oData <= 16'h0000;
            14'h1950: oData <= 16'ha000;
            14'h1951: oData <= 16'h02aa;
            14'h1952: oData <= 16'haa00;
            14'h1953: oData <= 16'h2a80;
            14'h1954: oData <= 16'h2aa0;
            14'h1955: oData <= 16'h0000;
            14'h1956: oData <= 16'h0000;
            14'h1957: oData <= 16'h0000;
            14'h1958: oData <= 16'h0000;
            14'h1959: oData <= 16'h0000;
            14'h195a: oData <= 16'haaa0;
            14'h195b: oData <= 16'h2aaa;
            14'h195c: oData <= 16'h0000;
            14'h195d: oData <= 16'h0000;
            14'h195e: oData <= 16'h0000;
            14'h195f: oData <= 16'h0000;
            14'h1960: oData <= 16'h0000;
            14'h1961: oData <= 16'h0000;
            14'h1962: oData <= 16'h0000;
            14'h1963: oData <= 16'h0000;
            14'h1964: oData <= 16'h8000;
            14'h1965: oData <= 16'h0aaa;
            14'h1966: oData <= 16'haa80;
            14'h1967: oData <= 16'h2aa0;
            14'h1968: oData <= 16'h0aa8;
            14'h1969: oData <= 16'h0000;
            14'h196a: oData <= 16'h0000;
            14'h196b: oData <= 16'h0000;
            14'h196c: oData <= 16'h0000;
            14'h196d: oData <= 16'ha800;
            14'h196e: oData <= 16'haaaa;
            14'h196f: oData <= 16'h0aaa;
            14'h1970: oData <= 16'h0000;
            14'h1971: oData <= 16'h0000;
            14'h1972: oData <= 16'h0000;
            14'h1973: oData <= 16'h0000;
            14'h1974: oData <= 16'h0000;
            14'h1975: oData <= 16'h0000;
            14'h1976: oData <= 16'h0000;
            14'h1977: oData <= 16'h0000;
            14'h1978: oData <= 16'h0000;
            14'h1979: oData <= 16'h0aaa;
            14'h197a: oData <= 16'haa80;
            14'h197b: oData <= 16'h2aa0;
            14'h197c: oData <= 16'h0aa8;
            14'h197d: oData <= 16'h0000;
            14'h197e: oData <= 16'h0000;
            14'h197f: oData <= 16'h0000;
            14'h1980: oData <= 16'h0000;
            14'h1981: oData <= 16'haaaa;
            14'h1982: oData <= 16'haaaa;
            14'h1983: oData <= 16'h02aa;
            14'h1984: oData <= 16'h0000;
            14'h1985: oData <= 16'h0000;
            14'h1986: oData <= 16'h0000;
            14'h1987: oData <= 16'h0000;
            14'h1988: oData <= 16'h0000;
            14'h1989: oData <= 16'h0000;
            14'h198a: oData <= 16'h0000;
            14'h198b: oData <= 16'h0000;
            14'h198c: oData <= 16'h0000;
            14'h198d: oData <= 16'haaa0;
            14'h198e: oData <= 16'h2a80;
            14'h198f: oData <= 16'h0aa8;
            14'h1990: oData <= 16'h02aa;
            14'h1991: oData <= 16'h0000;
            14'h1992: oData <= 16'h0000;
            14'h1993: oData <= 16'h0000;
            14'h1994: oData <= 16'haa80;
            14'h1995: oData <= 16'haaaa;
            14'h1996: oData <= 16'haaaa;
            14'h1997: oData <= 16'h00aa;
            14'h1998: oData <= 16'h0000;
            14'h1999: oData <= 16'h0000;
            14'h199a: oData <= 16'h0000;
            14'h199b: oData <= 16'h0000;
            14'h199c: oData <= 16'h0000;
            14'h199d: oData <= 16'h0000;
            14'h199e: oData <= 16'h0000;
            14'h199f: oData <= 16'h0000;
            14'h19a0: oData <= 16'h0000;
            14'h19a1: oData <= 16'haaa0;
            14'h19a2: oData <= 16'haa82;
            14'h19a3: oData <= 16'h0aaa;
            14'h19a4: oData <= 16'h02aa;
            14'h19a5: oData <= 16'h0000;
            14'h19a6: oData <= 16'h0000;
            14'h19a7: oData <= 16'ha000;
            14'h19a8: oData <= 16'haaaa;
            14'h19a9: oData <= 16'haaaa;
            14'h19aa: oData <= 16'haaaa;
            14'h19ab: oData <= 16'h00aa;
            14'h19ac: oData <= 16'h0000;
            14'h19ad: oData <= 16'h0000;
            14'h19ae: oData <= 16'h0000;
            14'h19af: oData <= 16'h0000;
            14'h19b0: oData <= 16'h0000;
            14'h19b1: oData <= 16'h0000;
            14'h19b2: oData <= 16'h0000;
            14'h19b3: oData <= 16'h0000;
            14'h19b4: oData <= 16'h0000;
            14'h19b5: oData <= 16'haa80;
            14'h19b6: oData <= 16'haa82;
            14'h19b7: oData <= 16'h0aaa;
            14'h19b8: oData <= 16'h00aa;
            14'h19b9: oData <= 16'h0000;
            14'h19ba: oData <= 16'ha000;
            14'h19bb: oData <= 16'haaaa;
            14'h19bc: oData <= 16'haaaa;
            14'h19bd: oData <= 16'haaaa;
            14'h19be: oData <= 16'h802a;
            14'h19bf: oData <= 16'h00aa;
            14'h19c0: oData <= 16'h0000;
            14'h19c1: oData <= 16'h0000;
            14'h19c2: oData <= 16'ha800;
            14'h19c3: oData <= 16'h0000;
            14'h19c4: oData <= 16'h0000;
            14'h19c5: oData <= 16'h0000;
            14'h19c6: oData <= 16'h0000;
            14'h19c7: oData <= 16'h0000;
            14'h19c8: oData <= 16'h0000;
            14'h19c9: oData <= 16'haa00;
            14'h19ca: oData <= 16'haa80;
            14'h19cb: oData <= 16'h82aa;
            14'h19cc: oData <= 16'h00aa;
            14'h19cd: oData <= 16'h0000;
            14'h19ce: oData <= 16'haa00;
            14'h19cf: oData <= 16'haaaa;
            14'h19d0: oData <= 16'haaaa;
            14'h19d1: oData <= 16'h0aaa;
            14'h19d2: oData <= 16'h8000;
            14'h19d3: oData <= 16'h00aa;
            14'h19d4: oData <= 16'h0000;
            14'h19d5: oData <= 16'h0000;
            14'h19d6: oData <= 16'haa80;
            14'h19d7: oData <= 16'h0002;
            14'h19d8: oData <= 16'h0000;
            14'h19d9: oData <= 16'h0000;
            14'h19da: oData <= 16'h0000;
            14'h19db: oData <= 16'h0000;
            14'h19dc: oData <= 16'h0000;
            14'h19dd: oData <= 16'h0000;
            14'h19de: oData <= 16'haa00;
            14'h19df: oData <= 16'h802a;
            14'h19e0: oData <= 16'h00aa;
            14'h19e1: oData <= 16'h0000;
            14'h19e2: oData <= 16'haaa0;
            14'h19e3: oData <= 16'haaaa;
            14'h19e4: oData <= 16'haaaa;
            14'h19e5: oData <= 16'h0002;
            14'h19e6: oData <= 16'h8000;
            14'h19e7: oData <= 16'h00aa;
            14'h19e8: oData <= 16'h0000;
            14'h19e9: oData <= 16'h0000;
            14'h19ea: oData <= 16'haaa8;
            14'h19eb: oData <= 16'h0002;
            14'h19ec: oData <= 16'h0000;
            14'h19ed: oData <= 16'h0000;
            14'h19ee: oData <= 16'h0000;
            14'h19ef: oData <= 16'h0000;
            14'h19f0: oData <= 16'h0000;
            14'h19f1: oData <= 16'h0000;
            14'h19f2: oData <= 16'ha000;
            14'h19f3: oData <= 16'h8002;
            14'h19f4: oData <= 16'h002a;
            14'h19f5: oData <= 16'h8000;
            14'h19f6: oData <= 16'haaaa;
            14'h19f7: oData <= 16'haaaa;
            14'h19f8: oData <= 16'h00aa;
            14'h19f9: oData <= 16'h0000;
            14'h19fa: oData <= 16'h8000;
            14'h19fb: oData <= 16'h02aa;
            14'h19fc: oData <= 16'h0000;
            14'h19fd: oData <= 16'h8000;
            14'h19fe: oData <= 16'haaaa;
            14'h19ff: oData <= 16'h000a;
            14'h1a00: oData <= 16'h0000;
            14'h1a01: oData <= 16'h0000;
            14'h1a02: oData <= 16'h0000;
            14'h1a03: oData <= 16'h0000;
            14'h1a04: oData <= 16'h0000;
            14'h1a05: oData <= 16'h0000;
            14'h1a06: oData <= 16'h0000;
            14'h1a07: oData <= 16'ha000;
            14'h1a08: oData <= 16'h002a;
            14'h1a09: oData <= 16'ha800;
            14'h1a0a: oData <= 16'haaaa;
            14'h1a0b: oData <= 16'h2aaa;
            14'h1a0c: oData <= 16'h0000;
            14'h1a0d: oData <= 16'h0000;
            14'h1a0e: oData <= 16'h0000;
            14'h1a0f: oData <= 16'h02aa;
            14'h1a10: oData <= 16'h0000;
            14'h1a11: oData <= 16'haa00;
            14'h1a12: oData <= 16'haaaa;
            14'h1a13: oData <= 16'h00aa;
            14'h1a14: oData <= 16'h0000;
            14'h1a15: oData <= 16'h0000;
            14'h1a16: oData <= 16'h0000;
            14'h1a17: oData <= 16'h0000;
            14'h1a18: oData <= 16'h0000;
            14'h1a19: oData <= 16'h0000;
            14'h1a1a: oData <= 16'h0000;
            14'h1a1b: oData <= 16'ha000;
            14'h1a1c: oData <= 16'h002a;
            14'h1a1d: oData <= 16'haaa0;
            14'h1a1e: oData <= 16'haaaa;
            14'h1a1f: oData <= 16'h0000;
            14'h1a20: oData <= 16'h0000;
            14'h1a21: oData <= 16'h0000;
            14'h1a22: oData <= 16'h0000;
            14'h1a23: oData <= 16'h02aa;
            14'h1a24: oData <= 16'h0000;
            14'h1a25: oData <= 16'haaa0;
            14'h1a26: oData <= 16'haaaa;
            14'h1a27: oData <= 16'h02aa;
            14'h1a28: oData <= 16'h0000;
            14'h1a29: oData <= 16'h0000;
            14'h1a2a: oData <= 16'h0000;
            14'h1a2b: oData <= 16'h0000;
            14'h1a2c: oData <= 16'h0000;
            14'h1a2d: oData <= 16'h0000;
            14'h1a2e: oData <= 16'h0000;
            14'h1a2f: oData <= 16'ha000;
            14'h1a30: oData <= 16'h000a;
            14'h1a31: oData <= 16'haaaa;
            14'h1a32: oData <= 16'h02aa;
            14'h1a33: oData <= 16'h0000;
            14'h1a34: oData <= 16'h0000;
            14'h1a35: oData <= 16'h0000;
            14'h1a36: oData <= 16'h0000;
            14'h1a37: oData <= 16'h02aa;
            14'h1a38: oData <= 16'h0000;
            14'h1a39: oData <= 16'haaaa;
            14'h1a3a: oData <= 16'h80aa;
            14'h1a3b: oData <= 16'h0aaa;
            14'h1a3c: oData <= 16'h0000;
            14'h1a3d: oData <= 16'h0000;
            14'h1a3e: oData <= 16'h0000;
            14'h1a3f: oData <= 16'h0000;
            14'h1a40: oData <= 16'h0000;
            14'h1a41: oData <= 16'h0000;
            14'h1a42: oData <= 16'h0000;
            14'h1a43: oData <= 16'ha800;
            14'h1a44: oData <= 16'ha80a;
            14'h1a45: oData <= 16'haaaa;
            14'h1a46: oData <= 16'h002a;
            14'h1a47: oData <= 16'h0000;
            14'h1a48: oData <= 16'h0000;
            14'h1a49: oData <= 16'h0000;
            14'h1a4a: oData <= 16'h0000;
            14'h1a4b: oData <= 16'h0aaa;
            14'h1a4c: oData <= 16'ha000;
            14'h1a4d: oData <= 16'haaaa;
            14'h1a4e: oData <= 16'h000a;
            14'h1a4f: oData <= 16'h2aaa;
            14'h1a50: oData <= 16'h0000;
            14'h1a51: oData <= 16'h0000;
            14'h1a52: oData <= 16'h0000;
            14'h1a53: oData <= 16'h0000;
            14'h1a54: oData <= 16'h0000;
            14'h1a55: oData <= 16'h0000;
            14'h1a56: oData <= 16'h0000;
            14'h1a57: oData <= 16'ha800;
            14'h1a58: oData <= 16'haaaa;
            14'h1a59: oData <= 16'haaaa;
            14'h1a5a: oData <= 16'h0000;
            14'h1a5b: oData <= 16'h0000;
            14'h1a5c: oData <= 16'h0000;
            14'h1a5d: oData <= 16'h0000;
            14'h1a5e: oData <= 16'h0000;
            14'h1a5f: oData <= 16'h0aa8;
            14'h1a60: oData <= 16'haa80;
            14'h1a61: oData <= 16'haaaa;
            14'h1a62: oData <= 16'h0000;
            14'h1a63: oData <= 16'haaa8;
            14'h1a64: oData <= 16'h0002;
            14'h1a65: oData <= 16'h0000;
            14'h1a66: oData <= 16'h0000;
            14'h1a67: oData <= 16'h0000;
            14'h1a68: oData <= 16'h0000;
            14'h1a69: oData <= 16'h0000;
            14'h1a6a: oData <= 16'h0000;
            14'h1a6b: oData <= 16'ha800;
            14'h1a6c: oData <= 16'haaaa;
            14'h1a6d: oData <= 16'h0aaa;
            14'h1a6e: oData <= 16'h0000;
            14'h1a6f: oData <= 16'h0000;
            14'h1a70: oData <= 16'h0000;
            14'h1a71: oData <= 16'h0000;
            14'h1a72: oData <= 16'h0000;
            14'h1a73: oData <= 16'h0aa8;
            14'h1a74: oData <= 16'haaa8;
            14'h1a75: oData <= 16'h02aa;
            14'h1a76: oData <= 16'h0000;
            14'h1a77: oData <= 16'haa80;
            14'h1a78: oData <= 16'h000a;
            14'h1a79: oData <= 16'h0000;
            14'h1a7a: oData <= 16'h0000;
            14'h1a7b: oData <= 16'h0000;
            14'h1a7c: oData <= 16'h0000;
            14'h1a7d: oData <= 16'h0000;
            14'h1a7e: oData <= 16'h0000;
            14'h1a7f: oData <= 16'ha800;
            14'h1a80: oData <= 16'haaaa;
            14'h1a81: oData <= 16'h002a;
            14'h1a82: oData <= 16'h0000;
            14'h1a83: oData <= 16'h0000;
            14'h1a84: oData <= 16'h0000;
            14'h1a85: oData <= 16'h0000;
            14'h1a86: oData <= 16'h0000;
            14'h1a87: oData <= 16'h8aa8;
            14'h1a88: oData <= 16'haaaa;
            14'h1a89: oData <= 16'h002a;
            14'h1a8a: oData <= 16'h0000;
            14'h1a8b: oData <= 16'haa00;
            14'h1a8c: oData <= 16'h002a;
            14'h1a8d: oData <= 16'h0000;
            14'h1a8e: oData <= 16'h0000;
            14'h1a8f: oData <= 16'h0000;
            14'h1a90: oData <= 16'h0000;
            14'h1a91: oData <= 16'h0000;
            14'h1a92: oData <= 16'h0000;
            14'h1a93: oData <= 16'ha800;
            14'h1a94: oData <= 16'haaaa;
            14'h1a95: oData <= 16'h0002;
            14'h1a96: oData <= 16'h0000;
            14'h1a97: oData <= 16'h0000;
            14'h1a98: oData <= 16'h0000;
            14'h1a99: oData <= 16'h0000;
            14'h1a9a: oData <= 16'h0000;
            14'h1a9b: oData <= 16'haaa8;
            14'h1a9c: oData <= 16'haaaa;
            14'h1a9d: oData <= 16'h0002;
            14'h1a9e: oData <= 16'h0000;
            14'h1a9f: oData <= 16'ha800;
            14'h1aa0: oData <= 16'h00aa;
            14'h1aa1: oData <= 16'h0000;
            14'h1aa2: oData <= 16'h0000;
            14'h1aa3: oData <= 16'h0000;
            14'h1aa4: oData <= 16'h0000;
            14'h1aa5: oData <= 16'h0000;
            14'h1aa6: oData <= 16'h0000;
            14'h1aa7: oData <= 16'ha800;
            14'h1aa8: oData <= 16'h0aaa;
            14'h1aa9: oData <= 16'h0000;
            14'h1aaa: oData <= 16'h0000;
            14'h1aab: oData <= 16'h0000;
            14'h1aac: oData <= 16'h0000;
            14'h1aad: oData <= 16'h0000;
            14'h1aae: oData <= 16'h0000;
            14'h1aaf: oData <= 16'haaa0;
            14'h1ab0: oData <= 16'h2aaa;
            14'h1ab1: oData <= 16'h0000;
            14'h1ab2: oData <= 16'h0000;
            14'h1ab3: oData <= 16'ha000;
            14'h1ab4: oData <= 16'h0aaa;
            14'h1ab5: oData <= 16'h0000;
            14'h1ab6: oData <= 16'h0000;
            14'h1ab7: oData <= 16'h0000;
            14'h1ab8: oData <= 16'h0000;
            14'h1ab9: oData <= 16'h0000;
            14'h1aba: oData <= 16'h0000;
            14'h1abb: oData <= 16'h8000;
            14'h1abc: oData <= 16'haaaa;
            14'h1abd: oData <= 16'h0000;
            14'h1abe: oData <= 16'h0000;
            14'h1abf: oData <= 16'h0000;
            14'h1ac0: oData <= 16'h0000;
            14'h1ac1: oData <= 16'h0000;
            14'h1ac2: oData <= 16'h0000;
            14'h1ac3: oData <= 16'haaa0;
            14'h1ac4: oData <= 16'h00aa;
            14'h1ac5: oData <= 16'h0000;
            14'h1ac6: oData <= 16'h0000;
            14'h1ac7: oData <= 16'h0000;
            14'h1ac8: oData <= 16'h2aaa;
            14'h1ac9: oData <= 16'h0000;
            14'h1aca: oData <= 16'h0000;
            14'h1acb: oData <= 16'h0000;
            14'h1acc: oData <= 16'h0000;
            14'h1acd: oData <= 16'h0000;
            14'h1ace: oData <= 16'h0000;
            14'h1acf: oData <= 16'h0000;
            14'h1ad0: oData <= 16'haaaa;
            14'h1ad1: oData <= 16'h0002;
            14'h1ad2: oData <= 16'h8000;
            14'h1ad3: oData <= 16'h000a;
            14'h1ad4: oData <= 16'h0000;
            14'h1ad5: oData <= 16'h0000;
            14'h1ad6: oData <= 16'h0000;
            14'h1ad7: oData <= 16'haaa0;
            14'h1ad8: oData <= 16'h000a;
            14'h1ad9: oData <= 16'h0000;
            14'h1ada: oData <= 16'h0000;
            14'h1adb: oData <= 16'h0000;
            14'h1adc: oData <= 16'haaa8;
            14'h1add: oData <= 16'h0000;
            14'h1ade: oData <= 16'h0000;
            14'h1adf: oData <= 16'h0000;
            14'h1ae0: oData <= 16'h0000;
            14'h1ae1: oData <= 16'h0000;
            14'h1ae2: oData <= 16'h0000;
            14'h1ae3: oData <= 16'h0000;
            14'h1ae4: oData <= 16'haaa0;
            14'h1ae5: oData <= 16'h0002;
            14'h1ae6: oData <= 16'ha000;
            14'h1ae7: oData <= 16'h002a;
            14'h1ae8: oData <= 16'h0000;
            14'h1ae9: oData <= 16'h0000;
            14'h1aea: oData <= 16'h0000;
            14'h1aeb: oData <= 16'haaaa;
            14'h1aec: oData <= 16'h0000;
            14'h1aed: oData <= 16'h0000;
            14'h1aee: oData <= 16'h0000;
            14'h1aef: oData <= 16'h0000;
            14'h1af0: oData <= 16'haaa0;
            14'h1af1: oData <= 16'h002a;
            14'h1af2: oData <= 16'h0000;
            14'h1af3: oData <= 16'h0000;
            14'h1af4: oData <= 16'h0000;
            14'h1af5: oData <= 16'h0000;
            14'h1af6: oData <= 16'h0000;
            14'h1af7: oData <= 16'h0000;
            14'h1af8: oData <= 16'haa00;
            14'h1af9: oData <= 16'h0000;
            14'h1afa: oData <= 16'ha000;
            14'h1afb: oData <= 16'h00aa;
            14'h1afc: oData <= 16'h0000;
            14'h1afd: oData <= 16'h0000;
            14'h1afe: oData <= 16'h8000;
            14'h1aff: oData <= 16'h2aaa;
            14'h1b00: oData <= 16'h0000;
            14'h1b01: oData <= 16'h0000;
            14'h1b02: oData <= 16'h0000;
            14'h1b03: oData <= 16'h0000;
            14'h1b04: oData <= 16'haa80;
            14'h1b05: oData <= 16'h00aa;
            14'h1b06: oData <= 16'h0000;
            14'h1b07: oData <= 16'h0000;
            14'h1b08: oData <= 16'h0000;
            14'h1b09: oData <= 16'h0000;
            14'h1b0a: oData <= 16'h0000;
            14'h1b0b: oData <= 16'h0000;
            14'h1b0c: oData <= 16'h0000;
            14'h1b0d: oData <= 16'h0000;
            14'h1b0e: oData <= 16'ha000;
            14'h1b0f: oData <= 16'h02aa;
            14'h1b10: oData <= 16'h0000;
            14'h1b11: oData <= 16'h0000;
            14'h1b12: oData <= 16'ha000;
            14'h1b13: oData <= 16'h0aaa;
            14'h1b14: oData <= 16'h0000;
            14'h1b15: oData <= 16'h0000;
            14'h1b16: oData <= 16'h0000;
            14'h1b17: oData <= 16'h0000;
            14'h1b18: oData <= 16'ha800;
            14'h1b19: oData <= 16'h00aa;
            14'h1b1a: oData <= 16'h0000;
            14'h1b1b: oData <= 16'h0000;
            14'h1b1c: oData <= 16'h0000;
            14'h1b1d: oData <= 16'h0000;
            14'h1b1e: oData <= 16'h0000;
            14'h1b1f: oData <= 16'h0000;
            14'h1b20: oData <= 16'h0000;
            14'h1b21: oData <= 16'h0000;
            14'h1b22: oData <= 16'h8000;
            14'h1b23: oData <= 16'h2aaa;
            14'h1b24: oData <= 16'h0000;
            14'h1b25: oData <= 16'h0000;
            14'h1b26: oData <= 16'haa00;
            14'h1b27: oData <= 16'h00aa;
            14'h1b28: oData <= 16'h0000;
            14'h1b29: oData <= 16'h0000;
            14'h1b2a: oData <= 16'h0000;
            14'h1b2b: oData <= 16'h0000;
            14'h1b2c: oData <= 16'ha000;
            14'h1b2d: oData <= 16'h00aa;
            14'h1b2e: oData <= 16'h0000;
            14'h1b2f: oData <= 16'h0000;
            14'h1b30: oData <= 16'h0000;
            14'h1b31: oData <= 16'h0000;
            14'h1b32: oData <= 16'h0000;
            14'h1b33: oData <= 16'h0000;
            14'h1b34: oData <= 16'h0000;
            14'h1b35: oData <= 16'h0000;
            14'h1b36: oData <= 16'h0000;
            14'h1b37: oData <= 16'haaaa;
            14'h1b38: oData <= 16'h0000;
            14'h1b39: oData <= 16'h0000;
            14'h1b3a: oData <= 16'haa80;
            14'h1b3b: oData <= 16'h002a;
            14'h1b3c: oData <= 16'h0000;
            14'h1b3d: oData <= 16'h0000;
            14'h1b3e: oData <= 16'h0000;
            14'h1b3f: oData <= 16'h0000;
            14'h1b40: oData <= 16'h8000;
            14'h1b41: oData <= 16'h002a;
            14'h1b42: oData <= 16'h0000;
            14'h1b43: oData <= 16'h0000;
            14'h1b44: oData <= 16'h0000;
            14'h1b45: oData <= 16'h0000;
            14'h1b46: oData <= 16'h0000;
            14'h1b47: oData <= 16'h0000;
            14'h1b48: oData <= 16'h0000;
            14'h1b49: oData <= 16'h0000;
            14'h1b4a: oData <= 16'h0000;
            14'h1b4b: oData <= 16'haaa8;
            14'h1b4c: oData <= 16'h000a;
            14'h1b4d: oData <= 16'h0000;
            14'h1b4e: oData <= 16'haaa0;
            14'h1b4f: oData <= 16'h0002;
            14'h1b50: oData <= 16'h0000;
            14'h1b51: oData <= 16'h0000;
            14'h1b52: oData <= 16'h0000;
            14'h1b53: oData <= 16'h0000;
            14'h1b54: oData <= 16'h0000;
            14'h1b55: oData <= 16'h0000;
            14'h1b56: oData <= 16'h0000;
            14'h1b57: oData <= 16'h0000;
            14'h1b58: oData <= 16'h0000;
            14'h1b59: oData <= 16'h0000;
            14'h1b5a: oData <= 16'h0000;
            14'h1b5b: oData <= 16'h0000;
            14'h1b5c: oData <= 16'h0000;
            14'h1b5d: oData <= 16'h0000;
            14'h1b5e: oData <= 16'h0000;
            14'h1b5f: oData <= 16'haa80;
            14'h1b60: oData <= 16'h002a;
            14'h1b61: oData <= 16'h0000;
            14'h1b62: oData <= 16'haaaa;
            14'h1b63: oData <= 16'h0000;
            14'h1b64: oData <= 16'h0000;
            14'h1b65: oData <= 16'h0000;
            14'h1b66: oData <= 16'h0000;
            14'h1b67: oData <= 16'h0000;
            14'h1b68: oData <= 16'h0000;
            14'h1b69: oData <= 16'h0000;
            14'h1b6a: oData <= 16'h0000;
            14'h1b6b: oData <= 16'h0000;
            14'h1b6c: oData <= 16'h0000;
            14'h1b6d: oData <= 16'h0000;
            14'h1b6e: oData <= 16'h0000;
            14'h1b6f: oData <= 16'h0000;
            14'h1b70: oData <= 16'h0000;
            14'h1b71: oData <= 16'h0000;
            14'h1b72: oData <= 16'h0000;
            14'h1b73: oData <= 16'haa00;
            14'h1b74: oData <= 16'h02aa;
            14'h1b75: oData <= 16'h8000;
            14'h1b76: oData <= 16'h2aaa;
            14'h1b77: oData <= 16'h0000;
            14'h1b78: oData <= 16'h0000;
            14'h1b79: oData <= 16'h0000;
            14'h1b7a: oData <= 16'h0000;
            14'h1b7b: oData <= 16'h0000;
            14'h1b7c: oData <= 16'h0000;
            14'h1b7d: oData <= 16'h0000;
            14'h1b7e: oData <= 16'h0000;
            14'h1b7f: oData <= 16'h0000;
            14'h1b80: oData <= 16'h0000;
            14'h1b81: oData <= 16'h0000;
            14'h1b82: oData <= 16'h0000;
            14'h1b83: oData <= 16'h0000;
            14'h1b84: oData <= 16'h0000;
            14'h1b85: oData <= 16'h0000;
            14'h1b86: oData <= 16'h0000;
            14'h1b87: oData <= 16'ha000;
            14'h1b88: oData <= 16'h0aaa;
            14'h1b89: oData <= 16'ha000;
            14'h1b8a: oData <= 16'h02aa;
            14'h1b8b: oData <= 16'h0000;
            14'h1b8c: oData <= 16'h0000;
            14'h1b8d: oData <= 16'h0000;
            14'h1b8e: oData <= 16'h0000;
            14'h1b8f: oData <= 16'h0000;
            14'h1b90: oData <= 16'h0000;
            14'h1b91: oData <= 16'h0000;
            14'h1b92: oData <= 16'h0000;
            14'h1b93: oData <= 16'h0000;
            14'h1b94: oData <= 16'h0000;
            14'h1b95: oData <= 16'h0000;
            14'h1b96: oData <= 16'h0000;
            14'h1b97: oData <= 16'h0000;
            14'h1b98: oData <= 16'h0000;
            14'h1b99: oData <= 16'h0000;
            14'h1b9a: oData <= 16'h0000;
            14'h1b9b: oData <= 16'h8000;
            14'h1b9c: oData <= 16'haaaa;
            14'h1b9d: oData <= 16'haa00;
            14'h1b9e: oData <= 16'h00aa;
            14'h1b9f: oData <= 16'h0000;
            14'h1ba0: oData <= 16'h0000;
            14'h1ba1: oData <= 16'h0000;
            14'h1ba2: oData <= 16'h0000;
            14'h1ba3: oData <= 16'h0000;
            14'h1ba4: oData <= 16'h0000;
            14'h1ba5: oData <= 16'h0000;
            14'h1ba6: oData <= 16'h0000;
            14'h1ba7: oData <= 16'h0000;
            14'h1ba8: oData <= 16'h0000;
            14'h1ba9: oData <= 16'h0000;
            14'h1baa: oData <= 16'h0000;
            14'h1bab: oData <= 16'h0000;
            14'h1bac: oData <= 16'h0000;
            14'h1bad: oData <= 16'h0000;
            14'h1bae: oData <= 16'h0000;
            14'h1baf: oData <= 16'h0000;
            14'h1bb0: oData <= 16'haaa8;
            14'h1bb1: oData <= 16'haa82;
            14'h1bb2: oData <= 16'h002a;
            14'h1bb3: oData <= 16'h0000;
            14'h1bb4: oData <= 16'h0000;
            14'h1bb5: oData <= 16'h0000;
            14'h1bb6: oData <= 16'h0000;
            14'h1bb7: oData <= 16'h0000;
            14'h1bb8: oData <= 16'h0000;
            14'h1bb9: oData <= 16'h0000;
            14'h1bba: oData <= 16'h0000;
            14'h1bbb: oData <= 16'h0000;
            14'h1bbc: oData <= 16'h0000;
            14'h1bbd: oData <= 16'h0000;
            14'h1bbe: oData <= 16'h0000;
            14'h1bbf: oData <= 16'h0000;
            14'h1bc0: oData <= 16'h0000;
            14'h1bc1: oData <= 16'h0000;
            14'h1bc2: oData <= 16'h0000;
            14'h1bc3: oData <= 16'h0000;
            14'h1bc4: oData <= 16'haaa0;
            14'h1bc5: oData <= 16'haaaa;
            14'h1bc6: oData <= 16'h0002;
            14'h1bc7: oData <= 16'h0000;
            14'h1bc8: oData <= 16'h0000;
            14'h1bc9: oData <= 16'h0000;
            14'h1bca: oData <= 16'h0000;
            14'h1bcb: oData <= 16'h0000;
            14'h1bcc: oData <= 16'h0000;
            14'h1bcd: oData <= 16'h0000;
            14'h1bce: oData <= 16'h0000;
            14'h1bcf: oData <= 16'h0000;
            14'h1bd0: oData <= 16'h0000;
            14'h1bd1: oData <= 16'h0000;
            14'h1bd2: oData <= 16'h0000;
            14'h1bd3: oData <= 16'h0000;
            14'h1bd4: oData <= 16'h0000;
            14'h1bd5: oData <= 16'h0000;
            14'h1bd6: oData <= 16'h0000;
            14'h1bd7: oData <= 16'h0000;
            14'h1bd8: oData <= 16'haa00;
            14'h1bd9: oData <= 16'haaaa;
            14'h1bda: oData <= 16'h0000;
            14'h1bdb: oData <= 16'h0000;
            14'h1bdc: oData <= 16'h0000;
            14'h1bdd: oData <= 16'h0000;
            14'h1bde: oData <= 16'h0000;
            14'h1bdf: oData <= 16'h0000;
            14'h1be0: oData <= 16'h0000;
            14'h1be1: oData <= 16'h0000;
            14'h1be2: oData <= 16'h0000;
            14'h1be3: oData <= 16'h0000;
            14'h1be4: oData <= 16'h0000;
            14'h1be5: oData <= 16'h0000;
            14'h1be6: oData <= 16'h0000;
            14'h1be7: oData <= 16'h0000;
            14'h1be8: oData <= 16'h0000;
            14'h1be9: oData <= 16'h0000;
            14'h1bea: oData <= 16'h0000;
            14'h1beb: oData <= 16'h0000;
            14'h1bec: oData <= 16'ha800;
            14'h1bed: oData <= 16'h2aaa;
            14'h1bee: oData <= 16'h0000;
            14'h1bef: oData <= 16'h0000;
            14'h1bf0: oData <= 16'h0000;
            14'h1bf1: oData <= 16'h0000;
            14'h1bf2: oData <= 16'h0000;
            14'h1bf3: oData <= 16'h0000;
            14'h1bf4: oData <= 16'h0000;
            14'h1bf5: oData <= 16'h0000;
            14'h1bf6: oData <= 16'h0000;
            14'h1bf7: oData <= 16'h0000;
            14'h1bf8: oData <= 16'h0000;
            14'h1bf9: oData <= 16'h0000;
            14'h1bfa: oData <= 16'h0000;
            14'h1bfb: oData <= 16'h0000;
            14'h1bfc: oData <= 16'h0000;
            14'h1bfd: oData <= 16'h0000;
            14'h1bfe: oData <= 16'h0000;
            14'h1bff: oData <= 16'h0000;
            14'h1c00: oData <= 16'h8000;
            14'h1c01: oData <= 16'h02aa;
            14'h1c02: oData <= 16'h0000;
            14'h1c03: oData <= 16'h0000;
            14'h1c04: oData <= 16'h0000;
            14'h1c05: oData <= 16'h0000;
            14'h1c06: oData <= 16'h0000;
            14'h1c07: oData <= 16'h0000;
            14'h1c08: oData <= 16'h0000;
            14'h1c09: oData <= 16'h0000;
            14'h1c0a: oData <= 16'h0000;
            14'h1c0b: oData <= 16'h0000;
            14'h1c0c: oData <= 16'h0000;
            14'h1c0d: oData <= 16'h0000;
            14'h1c0e: oData <= 16'h0000;
            14'h1c0f: oData <= 16'h0000;
            14'h1c10: oData <= 16'h0000;
            14'h1c11: oData <= 16'h0000;
            14'h1c12: oData <= 16'h0000;
            14'h1c13: oData <= 16'h0000;
            14'h1c14: oData <= 16'h0000;
            14'h1c15: oData <= 16'h00aa;
            14'h1c16: oData <= 16'h0000;
            14'h1c17: oData <= 16'h0000;
            14'h1c18: oData <= 16'h0000;
            14'h1c19: oData <= 16'h0000;
            14'h1c1a: oData <= 16'h0000;
            14'h1c1b: oData <= 16'h0000;
            14'h1c1c: oData <= 16'h0000;
            14'h1c1d: oData <= 16'h0000;
            14'h1c1e: oData <= 16'h0000;
            14'h1c1f: oData <= 16'h0000;
            14'h1c20: oData <= 16'h0000;
            14'h1c21: oData <= 16'h0000;
            14'h1c22: oData <= 16'h0000;
            14'h1c23: oData <= 16'h0000;
            14'h1c24: oData <= 16'h0000;
            14'h1c25: oData <= 16'h0000;
            14'h1c26: oData <= 16'h0000;
            14'h1c27: oData <= 16'h0000;
            14'h1c28: oData <= 16'h0000;
            14'h1c29: oData <= 16'h0000;
            14'h1c2a: oData <= 16'h0000;
            14'h1c2b: oData <= 16'h0000;
            14'h1c2c: oData <= 16'h0000;
            14'h1c2d: oData <= 16'h0000;
            14'h1c2e: oData <= 16'h0000;
            14'h1c2f: oData <= 16'h0000;
            14'h1c30: oData <= 16'h0000;
            14'h1c31: oData <= 16'h0000;
            14'h1c32: oData <= 16'h0000;
            14'h1c33: oData <= 16'h000a;
            14'h1c34: oData <= 16'h0000;
            14'h1c35: oData <= 16'h0000;
            14'h1c36: oData <= 16'h0000;
            14'h1c37: oData <= 16'h0000;
            14'h1c38: oData <= 16'h0000;
            14'h1c39: oData <= 16'h0000;
            14'h1c3a: oData <= 16'haaa0;
            14'h1c3b: oData <= 16'haaaa;
            14'h1c3c: oData <= 16'haaaa;
            14'h1c3d: oData <= 16'haaaa;
            14'h1c3e: oData <= 16'h0aaa;
            14'h1c3f: oData <= 16'h0000;
            14'h1c40: oData <= 16'h0000;
            14'h1c41: oData <= 16'h0000;
            14'h1c42: oData <= 16'h0000;
            14'h1c43: oData <= 16'h0000;
            14'h1c44: oData <= 16'h0000;
            14'h1c45: oData <= 16'h0000;
            14'h1c46: oData <= 16'h8000;
            14'h1c47: oData <= 16'h002a;
            14'h1c48: oData <= 16'h0000;
            14'h1c49: oData <= 16'h0000;
            14'h1c4a: oData <= 16'h0000;
            14'h1c4b: oData <= 16'h0000;
            14'h1c4c: oData <= 16'h0000;
            14'h1c4d: oData <= 16'h0000;
            14'h1c4e: oData <= 16'haaaa;
            14'h1c4f: oData <= 16'haaaa;
            14'h1c50: oData <= 16'haaaa;
            14'h1c51: oData <= 16'haaaa;
            14'h1c52: oData <= 16'haaaa;
            14'h1c53: oData <= 16'haaaa;
            14'h1c54: oData <= 16'h0002;
            14'h1c55: oData <= 16'h0000;
            14'h1c56: oData <= 16'h0000;
            14'h1c57: oData <= 16'h0000;
            14'h1c58: oData <= 16'h0000;
            14'h1c59: oData <= 16'h0000;
            14'h1c5a: oData <= 16'h8000;
            14'h1c5b: oData <= 16'h002a;
            14'h1c5c: oData <= 16'h0000;
            14'h1c5d: oData <= 16'h0000;
            14'h1c5e: oData <= 16'h0000;
            14'h1c5f: oData <= 16'h0000;
            14'h1c60: oData <= 16'h0000;
            14'h1c61: oData <= 16'ha000;
            14'h1c62: oData <= 16'hffea;
            14'h1c63: oData <= 16'hffff;
            14'h1c64: oData <= 16'hffff;
            14'h1c65: oData <= 16'hffff;
            14'h1c66: oData <= 16'habff;
            14'h1c67: oData <= 16'haaaa;
            14'h1c68: oData <= 16'h02aa;
            14'h1c69: oData <= 16'h0000;
            14'h1c6a: oData <= 16'h0000;
            14'h1c6b: oData <= 16'h0000;
            14'h1c6c: oData <= 16'h0000;
            14'h1c6d: oData <= 16'haa80;
            14'h1c6e: oData <= 16'h802a;
            14'h1c6f: oData <= 16'h002a;
            14'h1c70: oData <= 16'h0000;
            14'h1c71: oData <= 16'h0000;
            14'h1c72: oData <= 16'h0000;
            14'h1c73: oData <= 16'h0000;
            14'h1c74: oData <= 16'h0000;
            14'h1c75: oData <= 16'ha800;
            14'h1c76: oData <= 16'hfffe;
            14'h1c77: oData <= 16'hffff;
            14'h1c78: oData <= 16'haaaa;
            14'h1c79: oData <= 16'haaaa;
            14'h1c7a: oData <= 16'hfffe;
            14'h1c7b: oData <= 16'hffff;
            14'h1c7c: oData <= 16'haaaa;
            14'h1c7d: oData <= 16'h000a;
            14'h1c7e: oData <= 16'h0000;
            14'h1c7f: oData <= 16'h0000;
            14'h1c80: oData <= 16'h0000;
            14'h1c81: oData <= 16'haaa0;
            14'h1c82: oData <= 16'h80aa;
            14'h1c83: oData <= 16'h002a;
            14'h1c84: oData <= 16'h0000;
            14'h1c85: oData <= 16'h0000;
            14'h1c86: oData <= 16'h0000;
            14'h1c87: oData <= 16'h0000;
            14'h1c88: oData <= 16'h0000;
            14'h1c89: oData <= 16'hea00;
            14'h1c8a: oData <= 16'hffff;
            14'h1c8b: oData <= 16'habff;
            14'h1c8c: oData <= 16'hffff;
            14'h1c8d: oData <= 16'hffff;
            14'h1c8e: oData <= 16'haaab;
            14'h1c8f: oData <= 16'haaaa;
            14'h1c90: oData <= 16'haafe;
            14'h1c91: oData <= 16'h00aa;
            14'h1c92: oData <= 16'h0000;
            14'h1c93: oData <= 16'h0000;
            14'h1c94: oData <= 16'h0000;
            14'h1c95: oData <= 16'haaa8;
            14'h1c96: oData <= 16'h82aa;
            14'h1c97: oData <= 16'h002a;
            14'h1c98: oData <= 16'h0000;
            14'h1c99: oData <= 16'h0000;
            14'h1c9a: oData <= 16'h0000;
            14'h1c9b: oData <= 16'h0000;
            14'h1c9c: oData <= 16'h0000;
            14'h1c9d: oData <= 16'hfa80;
            14'h1c9e: oData <= 16'hffff;
            14'h1c9f: oData <= 16'hfebf;
            14'h1ca0: oData <= 16'habff;
            14'h1ca1: oData <= 16'hffaa;
            14'h1ca2: oData <= 16'hffff;
            14'h1ca3: oData <= 16'hffff;
            14'h1ca4: oData <= 16'hffff;
            14'h1ca5: oData <= 16'h02ab;
            14'h1ca6: oData <= 16'h0000;
            14'h1ca7: oData <= 16'h0000;
            14'h1ca8: oData <= 16'h0000;
            14'h1ca9: oData <= 16'haaa8;
            14'h1caa: oData <= 16'h8aaa;
            14'h1cab: oData <= 16'h002a;
            14'h1cac: oData <= 16'h0000;
            14'h1cad: oData <= 16'h0000;
            14'h1cae: oData <= 16'h0000;
            14'h1caf: oData <= 16'h0000;
            14'h1cb0: oData <= 16'h0000;
            14'h1cb1: oData <= 16'hfe80;
            14'h1cb2: oData <= 16'hffff;
            14'h1cb3: oData <= 16'hffeb;
            14'h1cb4: oData <= 16'hfeaa;
            14'h1cb5: oData <= 16'haaff;
            14'h1cb6: oData <= 16'hffff;
            14'h1cb7: oData <= 16'hffff;
            14'h1cb8: oData <= 16'heaab;
            14'h1cb9: oData <= 16'h2abf;
            14'h1cba: oData <= 16'h0000;
            14'h1cbb: oData <= 16'h00a8;
            14'h1cbc: oData <= 16'h0000;
            14'h1cbd: oData <= 16'h02a8;
            14'h1cbe: oData <= 16'h8aa8;
            14'h1cbf: oData <= 16'h282a;
            14'h1cc0: oData <= 16'h0000;
            14'h1cc1: oData <= 16'h0000;
            14'h1cc2: oData <= 16'h0000;
            14'h1cc3: oData <= 16'h0000;
            14'h1cc4: oData <= 16'h0000;
            14'h1cc5: oData <= 16'hfea0;
            14'h1cc6: oData <= 16'hbfff;
            14'h1cc7: oData <= 16'habfe;
            14'h1cc8: oData <= 16'hffff;
            14'h1cc9: oData <= 16'hffff;
            14'h1cca: oData <= 16'haaaa;
            14'h1ccb: oData <= 16'haaaa;
            14'h1ccc: oData <= 16'hbffe;
            14'h1ccd: oData <= 16'haafe;
            14'h1cce: oData <= 16'h0002;
            14'h1ccf: oData <= 16'h02aa;
            14'h1cd0: oData <= 16'h0000;
            14'h1cd1: oData <= 16'h02a8;
            14'h1cd2: oData <= 16'h8aa0;
            14'h1cd3: oData <= 16'haa2a;
            14'h1cd4: oData <= 16'h0000;
            14'h1cd5: oData <= 16'h0000;
            14'h1cd6: oData <= 16'h0000;
            14'h1cd7: oData <= 16'h0000;
            14'h1cd8: oData <= 16'h0000;
            14'h1cd9: oData <= 16'hffa8;
            14'h1cda: oData <= 16'hebff;
            14'h1cdb: oData <= 16'hfebf;
            14'h1cdc: oData <= 16'haabf;
            14'h1cdd: oData <= 16'hfeaa;
            14'h1cde: oData <= 16'hffff;
            14'h1cdf: oData <= 16'hffff;
            14'h1ce0: oData <= 16'hffff;
            14'h1ce1: oData <= 16'haffe;
            14'h1ce2: oData <= 16'h000a;
            14'h1ce3: oData <= 16'h02aa;
            14'h1ce4: oData <= 16'h0000;
            14'h1ce5: oData <= 16'h02a8;
            14'h1ce6: oData <= 16'h8aa0;
            14'h1ce7: oData <= 16'haaaa;
            14'h1ce8: oData <= 16'h0000;
            14'h1ce9: oData <= 16'h0000;
            14'h1cea: oData <= 16'h0000;
            14'h1ceb: oData <= 16'h0000;
            14'h1cec: oData <= 16'h0000;
            14'h1ced: oData <= 16'hffea;
            14'h1cee: oData <= 16'hfeff;
            14'h1cef: oData <= 16'hbfeb;
            14'h1cf0: oData <= 16'hffea;
            14'h1cf1: oData <= 16'hfaff;
            14'h1cf2: oData <= 16'hffff;
            14'h1cf3: oData <= 16'hffff;
            14'h1cf4: oData <= 16'hfeaa;
            14'h1cf5: oData <= 16'hffff;
            14'h1cf6: oData <= 16'h002a;
            14'h1cf7: oData <= 16'h00aa;
            14'h1cf8: oData <= 16'h0000;
            14'h1cf9: oData <= 16'h02a8;
            14'h1cfa: oData <= 16'h8aa0;
            14'h1cfb: oData <= 16'haaaa;
            14'h1cfc: oData <= 16'h0000;
            14'h1cfd: oData <= 16'h0000;
            14'h1cfe: oData <= 16'h0000;
            14'h1cff: oData <= 16'h0000;
            14'h1d00: oData <= 16'h0000;
            14'h1d01: oData <= 16'hfffa;
            14'h1d02: oData <= 16'hbfaf;
            14'h1d03: oData <= 16'heafe;
            14'h1d04: oData <= 16'hffff;
            14'h1d05: oData <= 16'hffaf;
            14'h1d06: oData <= 16'hffff;
            14'h1d07: oData <= 16'haabf;
            14'h1d08: oData <= 16'hfaff;
            14'h1d09: oData <= 16'hffff;
            14'h1d0a: oData <= 16'h00ab;
            14'h1d0b: oData <= 16'h00aa;
            14'h1d0c: oData <= 16'h0000;
            14'h1d0d: oData <= 16'h02a8;
            14'h1d0e: oData <= 16'h8aa0;
            14'h1d0f: oData <= 16'h2aaa;
            14'h1d10: oData <= 16'h0000;
            14'h1d11: oData <= 16'h0000;
            14'h1d12: oData <= 16'h0000;
            14'h1d13: oData <= 16'h0000;
            14'h1d14: oData <= 16'h8000;
            14'h1d15: oData <= 16'hfffa;
            14'h1d16: oData <= 16'heffb;
            14'h1d17: oData <= 16'hffaf;
            14'h1d18: oData <= 16'hffff;
            14'h1d19: oData <= 16'hfebf;
            14'h1d1a: oData <= 16'hffff;
            14'h1d1b: oData <= 16'hffea;
            14'h1d1c: oData <= 16'hafff;
            14'h1d1d: oData <= 16'hffff;
            14'h1d1e: oData <= 16'h00af;
            14'h1d1f: oData <= 16'h02aa;
            14'h1d20: oData <= 16'h0000;
            14'h1d21: oData <= 16'h02a8;
            14'h1d22: oData <= 16'h8aa0;
            14'h1d23: oData <= 16'h02aa;
            14'h1d24: oData <= 16'h0000;
            14'h1d25: oData <= 16'h0000;
            14'h1d26: oData <= 16'h0000;
            14'h1d27: oData <= 16'h0000;
            14'h1d28: oData <= 16'h8000;
            14'h1d29: oData <= 16'hfffe;
            14'h1d2a: oData <= 16'hfbfe;
            14'h1d2b: oData <= 16'hfffb;
            14'h1d2c: oData <= 16'hffff;
            14'h1d2d: oData <= 16'hfeff;
            14'h1d2e: oData <= 16'hffff;
            14'h1d2f: oData <= 16'hfffe;
            14'h1d30: oData <= 16'hffff;
            14'h1d31: oData <= 16'hfffe;
            14'h1d32: oData <= 16'h00af;
            14'h1d33: oData <= 16'h02aa;
            14'h1d34: oData <= 16'h0000;
            14'h1d35: oData <= 16'h2aa8;
            14'h1d36: oData <= 16'h0aa8;
            14'h1d37: oData <= 16'h00aa;
            14'h1d38: oData <= 16'h0000;
            14'h1d39: oData <= 16'h0000;
            14'h1d3a: oData <= 16'h0000;
            14'h1d3b: oData <= 16'h0000;
            14'h1d3c: oData <= 16'h8000;
            14'h1d3d: oData <= 16'hfffe;
            14'h1d3e: oData <= 16'hfeff;
            14'h1d3f: oData <= 16'hfffe;
            14'h1d40: oData <= 16'hffff;
            14'h1d41: oData <= 16'hfaff;
            14'h1d42: oData <= 16'hffff;
            14'h1d43: oData <= 16'hffbf;
            14'h1d44: oData <= 16'hffff;
            14'h1d45: oData <= 16'hfffe;
            14'h1d46: oData <= 16'h00af;
            14'h1d47: oData <= 16'h02a8;
            14'h1d48: oData <= 16'h0000;
            14'h1d49: oData <= 16'haaa8;
            14'h1d4a: oData <= 16'h0aaa;
            14'h1d4b: oData <= 16'h0000;
            14'h1d4c: oData <= 16'h0000;
            14'h1d4d: oData <= 16'h0000;
            14'h1d4e: oData <= 16'h0000;
            14'h1d4f: oData <= 16'h0000;
            14'h1d50: oData <= 16'ha000;
            14'h1d51: oData <= 16'hfffe;
            14'h1d52: oData <= 16'hbfbf;
            14'h1d53: oData <= 16'hffff;
            14'h1d54: oData <= 16'hffff;
            14'h1d55: oData <= 16'hfbff;
            14'h1d56: oData <= 16'hffff;
            14'h1d57: oData <= 16'hffef;
            14'h1d58: oData <= 16'hffff;
            14'h1d59: oData <= 16'hfffb;
            14'h1d5a: oData <= 16'h00af;
            14'h1d5b: oData <= 16'h02a8;
            14'h1d5c: oData <= 16'h0000;
            14'h1d5d: oData <= 16'haaa0;
            14'h1d5e: oData <= 16'h02aa;
            14'h1d5f: oData <= 16'h0000;
            14'h1d60: oData <= 16'h0000;
            14'h1d61: oData <= 16'h0000;
            14'h1d62: oData <= 16'h0000;
            14'h1d63: oData <= 16'h0000;
            14'h1d64: oData <= 16'ha000;
            14'h1d65: oData <= 16'hffff;
            14'h1d66: oData <= 16'hefff;
            14'h1d67: oData <= 16'hbfff;
            14'h1d68: oData <= 16'hfaaa;
            14'h1d69: oData <= 16'hfbff;
            14'h1d6a: oData <= 16'hffff;
            14'h1d6b: oData <= 16'hfffb;
            14'h1d6c: oData <= 16'hffff;
            14'h1d6d: oData <= 16'hfffb;
            14'h1d6e: oData <= 16'h02af;
            14'h1d6f: oData <= 16'h0aa8;
            14'h1d70: oData <= 16'h0000;
            14'h1d71: oData <= 16'haa80;
            14'h1d72: oData <= 16'h02aa;
            14'h1d73: oData <= 16'h0000;
            14'h1d74: oData <= 16'h0000;
            14'h1d75: oData <= 16'h0000;
            14'h1d76: oData <= 16'h0000;
            14'h1d77: oData <= 16'h0000;
            14'h1d78: oData <= 16'ha800;
            14'h1d79: oData <= 16'hffff;
            14'h1d7a: oData <= 16'hffff;
            14'h1d7b: oData <= 16'haabf;
            14'h1d7c: oData <= 16'haaaa;
            14'h1d7d: oData <= 16'hfbfe;
            14'h1d7e: oData <= 16'hffff;
            14'h1d7f: oData <= 16'hfffb;
            14'h1d80: oData <= 16'hffff;
            14'h1d81: oData <= 16'hffff;
            14'h1d82: oData <= 16'h02bf;
            14'h1d83: oData <= 16'h0aa8;
            14'h1d84: oData <= 16'h0000;
            14'h1d85: oData <= 16'ha800;
            14'h1d86: oData <= 16'h002a;
            14'h1d87: oData <= 16'h0000;
            14'h1d88: oData <= 16'h0000;
            14'h1d89: oData <= 16'h0000;
            14'h1d8a: oData <= 16'h0000;
            14'h1d8b: oData <= 16'h0000;
            14'h1d8c: oData <= 16'hea00;
            14'h1d8d: oData <= 16'hffff;
            14'h1d8e: oData <= 16'hffff;
            14'h1d8f: oData <= 16'haaab;
            14'h1d90: oData <= 16'habaa;
            14'h1d91: oData <= 16'hffea;
            14'h1d92: oData <= 16'hffff;
            14'h1d93: oData <= 16'hfffb;
            14'h1d94: oData <= 16'hffff;
            14'h1d95: oData <= 16'hffff;
            14'h1d96: oData <= 16'h02bf;
            14'h1d97: oData <= 16'h2aa0;
            14'h1d98: oData <= 16'h0000;
            14'h1d99: oData <= 16'h0000;
            14'h1d9a: oData <= 16'h0000;
            14'h1d9b: oData <= 16'h0000;
            14'h1d9c: oData <= 16'h0000;
            14'h1d9d: oData <= 16'h0000;
            14'h1d9e: oData <= 16'h0000;
            14'h1d9f: oData <= 16'h0000;
            14'h1da0: oData <= 16'hfa80;
            14'h1da1: oData <= 16'hffff;
            14'h1da2: oData <= 16'hffff;
            14'h1da3: oData <= 16'haaaa;
            14'h1da4: oData <= 16'hffaa;
            14'h1da5: oData <= 16'hffaa;
            14'h1da6: oData <= 16'hffff;
            14'h1da7: oData <= 16'habfb;
            14'h1da8: oData <= 16'heaaa;
            14'h1da9: oData <= 16'hffff;
            14'h1daa: oData <= 16'h0abf;
            14'h1dab: oData <= 16'h2aa0;
            14'h1dac: oData <= 16'h0000;
            14'h1dad: oData <= 16'h0000;
            14'h1dae: oData <= 16'h0000;
            14'h1daf: oData <= 16'h0000;
            14'h1db0: oData <= 16'h0000;
            14'h1db1: oData <= 16'h0000;
            14'h1db2: oData <= 16'h0000;
            14'h1db3: oData <= 16'h0000;
            14'h1db4: oData <= 16'haaa0;
            14'h1db5: oData <= 16'hffea;
            14'h1db6: oData <= 16'hbebf;
            14'h1db7: oData <= 16'haafa;
            14'h1db8: oData <= 16'hffaa;
            14'h1db9: oData <= 16'hfaaf;
            14'h1dba: oData <= 16'hffff;
            14'h1dbb: oData <= 16'haabf;
            14'h1dbc: oData <= 16'haffe;
            14'h1dbd: oData <= 16'hfffe;
            14'h1dbe: oData <= 16'haaff;
            14'h1dbf: oData <= 16'haa80;
            14'h1dc0: oData <= 16'h0000;
            14'h1dc1: oData <= 16'h000a;
            14'h1dc2: oData <= 16'h0000;
            14'h1dc3: oData <= 16'h0000;
            14'h1dc4: oData <= 16'h0000;
            14'h1dc5: oData <= 16'h0000;
            14'h1dc6: oData <= 16'h0000;
            14'h1dc7: oData <= 16'h0000;
            14'h1dc8: oData <= 16'hfea8;
            14'h1dc9: oData <= 16'hffff;
            14'h1dca: oData <= 16'hafeb;
            14'h1dcb: oData <= 16'haaaa;
            14'h1dcc: oData <= 16'hfaaa;
            14'h1dcd: oData <= 16'hfabf;
            14'h1dce: oData <= 16'hffff;
            14'h1dcf: oData <= 16'haaaf;
            14'h1dd0: oData <= 16'haaaa;
            14'h1dd1: oData <= 16'hffbe;
            14'h1dd2: oData <= 16'habff;
            14'h1dd3: oData <= 16'haa82;
            14'h1dd4: oData <= 16'ha800;
            14'h1dd5: oData <= 16'h002a;
            14'h1dd6: oData <= 16'h0000;
            14'h1dd7: oData <= 16'h0000;
            14'h1dd8: oData <= 16'h0000;
            14'h1dd9: oData <= 16'h0000;
            14'h1dda: oData <= 16'h0000;
            14'h1ddb: oData <= 16'h0000;
            14'h1ddc: oData <= 16'haaea;
            14'h1ddd: oData <= 16'hfeaa;
            14'h1dde: oData <= 16'hafaf;
            14'h1ddf: oData <= 16'haaaa;
            14'h1de0: oData <= 16'haaaa;
            14'h1de1: oData <= 16'heaff;
            14'h1de2: oData <= 16'hafff;
            14'h1de3: oData <= 16'haaab;
            14'h1de4: oData <= 16'haaaa;
            14'h1de5: oData <= 16'haeae;
            14'h1de6: oData <= 16'hbfaa;
            14'h1de7: oData <= 16'haa0a;
            14'h1de8: oData <= 16'haa82;
            14'h1de9: oData <= 16'h002a;
            14'h1dea: oData <= 16'h0000;
            14'h1deb: oData <= 16'h0000;
            14'h1dec: oData <= 16'h0000;
            14'h1ded: oData <= 16'h0000;
            14'h1dee: oData <= 16'h0000;
            14'h1def: oData <= 16'h8000;
            14'h1df0: oData <= 16'hffba;
            14'h1df1: oData <= 16'hffff;
            14'h1df2: oData <= 16'hfaff;
            14'h1df3: oData <= 16'hfffa;
            14'h1df4: oData <= 16'habff;
            14'h1df5: oData <= 16'hfaaa;
            14'h1df6: oData <= 16'habff;
            14'h1df7: oData <= 16'haaaa;
            14'h1df8: oData <= 16'hfffa;
            14'h1df9: oData <= 16'hfbff;
            14'h1dfa: oData <= 16'hfeff;
            14'h1dfb: oData <= 16'haa0a;
            14'h1dfc: oData <= 16'haaaa;
            14'h1dfd: oData <= 16'h002a;
            14'h1dfe: oData <= 16'h0000;
            14'h1dff: oData <= 16'h0000;
            14'h1e00: oData <= 16'h0000;
            14'h1e01: oData <= 16'h0000;
            14'h1e02: oData <= 16'h0000;
            14'h1e03: oData <= 16'ha000;
            14'h1e04: oData <= 16'hffee;
            14'h1e05: oData <= 16'haaaa;
            14'h1e06: oData <= 16'hfeff;
            14'h1e07: oData <= 16'hbfff;
            14'h1e08: oData <= 16'hbffa;
            14'h1e09: oData <= 16'hfaaa;
            14'h1e0a: oData <= 16'hbfff;
            14'h1e0b: oData <= 16'hfeaa;
            14'h1e0c: oData <= 16'hffff;
            14'h1e0d: oData <= 16'hffff;
            14'h1e0e: oData <= 16'hfbeb;
            14'h1e0f: oData <= 16'ha82a;
            14'h1e10: oData <= 16'haaaa;
            14'h1e11: oData <= 16'h000a;
            14'h1e12: oData <= 16'h0000;
            14'h1e13: oData <= 16'h0000;
            14'h1e14: oData <= 16'h0000;
            14'h1e15: oData <= 16'h0000;
            14'h1e16: oData <= 16'h0000;
            14'h1e17: oData <= 16'ha800;
            14'h1e18: oData <= 16'haffb;
            14'h1e19: oData <= 16'haaaa;
            14'h1e1a: oData <= 16'hffea;
            14'h1e1b: oData <= 16'hafff;
            14'h1e1c: oData <= 16'hfffe;
            14'h1e1d: oData <= 16'hffaf;
            14'h1e1e: oData <= 16'hffff;
            14'h1e1f: oData <= 16'hffeb;
            14'h1e20: oData <= 16'hffff;
            14'h1e21: oData <= 16'hffff;
            14'h1e22: oData <= 16'hafbf;
            14'h1e23: oData <= 16'ha02b;
            14'h1e24: oData <= 16'h2aaa;
            14'h1e25: oData <= 16'h0000;
            14'h1e26: oData <= 16'h0000;
            14'h1e27: oData <= 16'h0000;
            14'h1e28: oData <= 16'h0000;
            14'h1e29: oData <= 16'h0000;
            14'h1e2a: oData <= 16'h0000;
            14'h1e2b: oData <= 16'he800;
            14'h1e2c: oData <= 16'habfe;
            14'h1e2d: oData <= 16'hbffe;
            14'h1e2e: oData <= 16'hfeaa;
            14'h1e2f: oData <= 16'haaff;
            14'h1e30: oData <= 16'hffff;
            14'h1e31: oData <= 16'hffff;
            14'h1e32: oData <= 16'hffff;
            14'h1e33: oData <= 16'hffeb;
            14'h1e34: oData <= 16'hffff;
            14'h1e35: oData <= 16'haabf;
            14'h1e36: oData <= 16'hbefe;
            14'h1e37: oData <= 16'h802b;
            14'h1e38: oData <= 16'h02aa;
            14'h1e39: oData <= 16'h0000;
            14'h1e3a: oData <= 16'h0000;
            14'h1e3b: oData <= 16'h0000;
            14'h1e3c: oData <= 16'h0000;
            14'h1e3d: oData <= 16'h0000;
            14'h1e3e: oData <= 16'h0000;
            14'h1e3f: oData <= 16'hea00;
            14'h1e40: oData <= 16'hebfe;
            14'h1e41: oData <= 16'hfbff;
            14'h1e42: oData <= 16'haaab;
            14'h1e43: oData <= 16'heaaa;
            14'h1e44: oData <= 16'hffff;
            14'h1e45: oData <= 16'hffff;
            14'h1e46: oData <= 16'hffff;
            14'h1e47: oData <= 16'hffeb;
            14'h1e48: oData <= 16'hffff;
            14'h1e49: oData <= 16'haaaf;
            14'h1e4a: oData <= 16'hfeea;
            14'h1e4b: oData <= 16'h002a;
            14'h1e4c: oData <= 16'h0000;
            14'h1e4d: oData <= 16'h0000;
            14'h1e4e: oData <= 16'h0000;
            14'h1e4f: oData <= 16'h0000;
            14'h1e50: oData <= 16'h0000;
            14'h1e51: oData <= 16'h0000;
            14'h1e52: oData <= 16'h0000;
            14'h1e53: oData <= 16'hfa00;
            14'h1e54: oData <= 16'heafe;
            14'h1e55: oData <= 16'hfaff;
            14'h1e56: oData <= 16'haaff;
            14'h1e57: oData <= 16'hfeaa;
            14'h1e58: oData <= 16'hffff;
            14'h1e59: oData <= 16'hffff;
            14'h1e5a: oData <= 16'hffff;
            14'h1e5b: oData <= 16'hffeb;
            14'h1e5c: oData <= 16'hfebf;
            14'h1e5d: oData <= 16'hffaa;
            14'h1e5e: oData <= 16'hfeea;
            14'h1e5f: oData <= 16'h002a;
            14'h1e60: oData <= 16'h0000;
            14'h1e61: oData <= 16'h0000;
            14'h1e62: oData <= 16'h0000;
            14'h1e63: oData <= 16'h0000;
            14'h1e64: oData <= 16'h0000;
            14'h1e65: oData <= 16'h0000;
            14'h1e66: oData <= 16'h0000;
            14'h1e67: oData <= 16'hfa80;
            14'h1e68: oData <= 16'hfafe;
            14'h1e69: oData <= 16'hfaff;
            14'h1e6a: oData <= 16'hffff;
            14'h1e6b: oData <= 16'hffff;
            14'h1e6c: oData <= 16'hffff;
            14'h1e6d: oData <= 16'hffff;
            14'h1e6e: oData <= 16'hffff;
            14'h1e6f: oData <= 16'hffeb;
            14'h1e70: oData <= 16'haabf;
            14'h1e71: oData <= 16'hffea;
            14'h1e72: oData <= 16'hfeef;
            14'h1e73: oData <= 16'h002a;
            14'h1e74: oData <= 16'h0000;
            14'h1e75: oData <= 16'h0000;
            14'h1e76: oData <= 16'h0000;
            14'h1e77: oData <= 16'h0000;
            14'h1e78: oData <= 16'h0000;
            14'h1e79: oData <= 16'h0000;
            14'h1e7a: oData <= 16'h0000;
            14'h1e7b: oData <= 16'hfe80;
            14'h1e7c: oData <= 16'hfabe;
            14'h1e7d: oData <= 16'haaff;
            14'h1e7e: oData <= 16'hffff;
            14'h1e7f: oData <= 16'hffff;
            14'h1e80: oData <= 16'hffff;
            14'h1e81: oData <= 16'hffff;
            14'h1e82: oData <= 16'hffff;
            14'h1e83: oData <= 16'hfeab;
            14'h1e84: oData <= 16'haaff;
            14'h1e85: oData <= 16'hfbfa;
            14'h1e86: oData <= 16'hfbff;
            14'h1e87: oData <= 16'h002a;
            14'h1e88: oData <= 16'h0000;
            14'h1e89: oData <= 16'h0000;
            14'h1e8a: oData <= 16'h0000;
            14'h1e8b: oData <= 16'h0000;
            14'h1e8c: oData <= 16'h0000;
            14'h1e8d: oData <= 16'h0000;
            14'h1e8e: oData <= 16'h0000;
            14'h1e8f: oData <= 16'hfe80;
            14'h1e90: oData <= 16'hfebe;
            14'h1e91: oData <= 16'haabf;
            14'h1e92: oData <= 16'hfffa;
            14'h1e93: oData <= 16'hffff;
            14'h1e94: oData <= 16'hefff;
            14'h1e95: oData <= 16'hfeab;
            14'h1e96: oData <= 16'hffff;
            14'h1e97: oData <= 16'hfaaf;
            14'h1e98: oData <= 16'hffff;
            14'h1e99: oData <= 16'hfaff;
            14'h1e9a: oData <= 16'hfbff;
            14'h1e9b: oData <= 16'h002a;
            14'h1e9c: oData <= 16'h0000;
            14'h1e9d: oData <= 16'h0000;
            14'h1e9e: oData <= 16'h0000;
            14'h1e9f: oData <= 16'h0000;
            14'h1ea0: oData <= 16'h0000;
            14'h1ea1: oData <= 16'h0000;
            14'h1ea2: oData <= 16'h0000;
            14'h1ea3: oData <= 16'hfe80;
            14'h1ea4: oData <= 16'hfebe;
            14'h1ea5: oData <= 16'hbeab;
            14'h1ea6: oData <= 16'hffaa;
            14'h1ea7: oData <= 16'hffff;
            14'h1ea8: oData <= 16'hefff;
            14'h1ea9: oData <= 16'hfaaa;
            14'h1eaa: oData <= 16'hffff;
            14'h1eab: oData <= 16'haaff;
            14'h1eac: oData <= 16'hffff;
            14'h1ead: oData <= 16'hfaff;
            14'h1eae: oData <= 16'hfbff;
            14'h1eaf: oData <= 16'h002a;
            14'h1eb0: oData <= 16'h0000;
            14'h1eb1: oData <= 16'h0000;
            14'h1eb2: oData <= 16'h0000;
            14'h1eb3: oData <= 16'h0000;
            14'h1eb4: oData <= 16'h0000;
            14'h1eb5: oData <= 16'h0000;
            14'h1eb6: oData <= 16'h0000;
            14'h1eb7: oData <= 16'hfa80;
            14'h1eb8: oData <= 16'hbebe;
            14'h1eb9: oData <= 16'hfeaa;
            14'h1eba: oData <= 16'hfaab;
            14'h1ebb: oData <= 16'hafff;
            14'h1ebc: oData <= 16'hbaaa;
            14'h1ebd: oData <= 16'hfffa;
            14'h1ebe: oData <= 16'hffff;
            14'h1ebf: oData <= 16'habff;
            14'h1ec0: oData <= 16'hfffe;
            14'h1ec1: oData <= 16'hfaff;
            14'h1ec2: oData <= 16'hbeff;
            14'h1ec3: oData <= 16'h002b;
            14'h1ec4: oData <= 16'h0000;
            14'h1ec5: oData <= 16'h0000;
            14'h1ec6: oData <= 16'h0000;
            14'h1ec7: oData <= 16'h0000;
            14'h1ec8: oData <= 16'h0000;
            14'h1ec9: oData <= 16'h0000;
            14'h1eca: oData <= 16'h0000;
            14'h1ecb: oData <= 16'hfa00;
            14'h1ecc: oData <= 16'hbabe;
            14'h1ecd: oData <= 16'hfaba;
            14'h1ece: oData <= 16'haabf;
            14'h1ecf: oData <= 16'heffe;
            14'h1ed0: oData <= 16'hbfff;
            14'h1ed1: oData <= 16'hfffe;
            14'h1ed2: oData <= 16'hffff;
            14'h1ed3: oData <= 16'habff;
            14'h1ed4: oData <= 16'hfffa;
            14'h1ed5: oData <= 16'haaff;
            14'h1ed6: oData <= 16'hbfaf;
            14'h1ed7: oData <= 16'h002a;
            14'h1ed8: oData <= 16'h0000;
            14'h1ed9: oData <= 16'h0000;
            14'h1eda: oData <= 16'h0000;
            14'h1edb: oData <= 16'h0000;
            14'h1edc: oData <= 16'h0000;
            14'h1edd: oData <= 16'h0000;
            14'h1ede: oData <= 16'h0000;
            14'h1edf: oData <= 16'hfa00;
            14'h1ee0: oData <= 16'hfafe;
            14'h1ee1: oData <= 16'hfaff;
            14'h1ee2: oData <= 16'habff;
            14'h1ee3: oData <= 16'hffea;
            14'h1ee4: oData <= 16'hbfff;
            14'h1ee5: oData <= 16'haafe;
            14'h1ee6: oData <= 16'hffea;
            14'h1ee7: oData <= 16'haaff;
            14'h1ee8: oData <= 16'hffae;
            14'h1ee9: oData <= 16'haaff;
            14'h1eea: oData <= 16'hefff;
            14'h1eeb: oData <= 16'h000a;
            14'h1eec: oData <= 16'h0000;
            14'h1eed: oData <= 16'h0000;
            14'h1eee: oData <= 16'h0000;
            14'h1eef: oData <= 16'h0000;
            14'h1ef0: oData <= 16'h0000;
            14'h1ef1: oData <= 16'h0000;
            14'h1ef2: oData <= 16'h0000;
            14'h1ef3: oData <= 16'hfa00;
            14'h1ef4: oData <= 16'heafb;
            14'h1ef5: oData <= 16'heaff;
            14'h1ef6: oData <= 16'hbfff;
            14'h1ef7: oData <= 16'hfaaa;
            14'h1ef8: oData <= 16'hbfff;
            14'h1ef9: oData <= 16'haafa;
            14'h1efa: oData <= 16'hffea;
            14'h1efb: oData <= 16'hbaff;
            14'h1efc: oData <= 16'hfafe;
            14'h1efd: oData <= 16'haabf;
            14'h1efe: oData <= 16'hfabf;
            14'h1eff: oData <= 16'h000a;
            14'h1f00: oData <= 16'h0000;
            14'h1f01: oData <= 16'h0000;
            14'h1f02: oData <= 16'h0000;
            14'h1f03: oData <= 16'h0000;
            14'h1f04: oData <= 16'h0000;
            14'h1f05: oData <= 16'h0000;
            14'h1f06: oData <= 16'h0000;
            14'h1f07: oData <= 16'hea00;
            14'h1f08: oData <= 16'hebfb;
            14'h1f09: oData <= 16'haaff;
            14'h1f0a: oData <= 16'hbfff;
            14'h1f0b: oData <= 16'haaae;
            14'h1f0c: oData <= 16'hfffa;
            14'h1f0d: oData <= 16'hfeea;
            14'h1f0e: oData <= 16'hffff;
            14'h1f0f: oData <= 16'hfabf;
            14'h1f10: oData <= 16'hefff;
            14'h1f11: oData <= 16'haeaf;
            14'h1f12: oData <= 16'hbfef;
            14'h1f13: oData <= 16'h000a;
            14'h1f14: oData <= 16'h0000;
            14'h1f15: oData <= 16'h0000;
            14'h1f16: oData <= 16'h0000;
            14'h1f17: oData <= 16'h0000;
            14'h1f18: oData <= 16'h0000;
            14'h1f19: oData <= 16'h0000;
            14'h1f1a: oData <= 16'h0000;
            14'h1f1b: oData <= 16'ha800;
            14'h1f1c: oData <= 16'hffef;
            14'h1f1d: oData <= 16'haaff;
            14'h1f1e: oData <= 16'hbffa;
            14'h1f1f: oData <= 16'habfe;
            14'h1f20: oData <= 16'hfeaa;
            14'h1f21: oData <= 16'hfffb;
            14'h1f22: oData <= 16'hafff;
            14'h1f23: oData <= 16'hfeab;
            14'h1f24: oData <= 16'hffff;
            14'h1f25: oData <= 16'haaab;
            14'h1f26: oData <= 16'hafff;
            14'h1f27: oData <= 16'h0002;
            14'h1f28: oData <= 16'h0000;
            14'h1f29: oData <= 16'h0000;
            14'h1f2a: oData <= 16'h0000;
            14'h1f2b: oData <= 16'h0000;
            14'h1f2c: oData <= 16'h0000;
            14'h1f2d: oData <= 16'h0000;
            14'h1f2e: oData <= 16'h0000;
            14'h1f2f: oData <= 16'ha000;
            14'h1f30: oData <= 16'hfebf;
            14'h1f31: oData <= 16'habff;
            14'h1f32: oData <= 16'hbfaa;
            14'h1f33: oData <= 16'hfffe;
            14'h1f34: oData <= 16'haaab;
            14'h1f35: oData <= 16'hffff;
            14'h1f36: oData <= 16'hafff;
            14'h1f37: oData <= 16'hffaa;
            14'h1f38: oData <= 16'hbfff;
            14'h1f39: oData <= 16'haaea;
            14'h1f3a: oData <= 16'haffe;
            14'h1f3b: oData <= 16'h0000;
            14'h1f3c: oData <= 16'h0000;
            14'h1f3d: oData <= 16'h0000;
            14'h1f3e: oData <= 16'h0000;
            14'h1f3f: oData <= 16'h0000;
            14'h1f40: oData <= 16'h0000;
            14'h1f41: oData <= 16'h0000;
            14'h1f42: oData <= 16'h0000;
            14'h1f43: oData <= 16'ha000;
            14'h1f44: oData <= 16'hebfe;
            14'h1f45: oData <= 16'hafff;
            14'h1f46: oData <= 16'hbaaa;
            14'h1f47: oData <= 16'hfffa;
            14'h1f48: oData <= 16'haaff;
            14'h1f49: oData <= 16'hffaa;
            14'h1f4a: oData <= 16'hbfff;
            14'h1f4b: oData <= 16'hfffa;
            14'h1f4c: oData <= 16'habff;
            14'h1f4d: oData <= 16'hbaea;
            14'h1f4e: oData <= 16'habfe;
            14'h1f4f: oData <= 16'h0000;
            14'h1f50: oData <= 16'h0000;
            14'h1f51: oData <= 16'h0000;
            14'h1f52: oData <= 16'h0000;
            14'h1f53: oData <= 16'h0000;
            14'h1f54: oData <= 16'h0000;
            14'h1f55: oData <= 16'h0000;
            14'h1f56: oData <= 16'h0000;
            14'h1f57: oData <= 16'h8000;
            14'h1f58: oData <= 16'hffaa;
            14'h1f59: oData <= 16'hbfff;
            14'h1f5a: oData <= 16'haaae;
            14'h1f5b: oData <= 16'hffea;
            14'h1f5c: oData <= 16'habff;
            14'h1f5d: oData <= 16'haaaa;
            14'h1f5e: oData <= 16'hfffa;
            14'h1f5f: oData <= 16'hffff;
            14'h1f60: oData <= 16'haaaf;
            14'h1f61: oData <= 16'haaeb;
            14'h1f62: oData <= 16'h2bfe;
            14'h1f63: oData <= 16'h0000;
            14'h1f64: oData <= 16'h0000;
            14'h1f65: oData <= 16'h0000;
            14'h1f66: oData <= 16'h0000;
            14'h1f67: oData <= 16'h0000;
            14'h1f68: oData <= 16'h0000;
            14'h1f69: oData <= 16'h0000;
            14'h1f6a: oData <= 16'h0000;
            14'h1f6b: oData <= 16'h0000;
            14'h1f6c: oData <= 16'hfeea;
            14'h1f6d: oData <= 16'hbfff;
            14'h1f6e: oData <= 16'habfa;
            14'h1f6f: oData <= 16'hffaa;
            14'h1f70: oData <= 16'hebff;
            14'h1f71: oData <= 16'haabf;
            14'h1f72: oData <= 16'haaaa;
            14'h1f73: oData <= 16'haaaa;
            14'h1f74: oData <= 16'hfaaa;
            14'h1f75: oData <= 16'habeb;
            14'h1f76: oData <= 16'h2bfe;
            14'h1f77: oData <= 16'h0000;
            14'h1f78: oData <= 16'h0000;
            14'h1f79: oData <= 16'h0000;
            14'h1f7a: oData <= 16'h0000;
            14'h1f7b: oData <= 16'h0000;
            14'h1f7c: oData <= 16'h0000;
            14'h1f7d: oData <= 16'h0000;
            14'h1f7e: oData <= 16'h0000;
            14'h1f7f: oData <= 16'h0000;
            14'h1f80: oData <= 16'hffa8;
            14'h1f81: oData <= 16'hffff;
            14'h1f82: oData <= 16'hbfea;
            14'h1f83: oData <= 16'heaaa;
            14'h1f84: oData <= 16'hebff;
            14'h1f85: oData <= 16'hffff;
            14'h1f86: oData <= 16'haaab;
            14'h1f87: oData <= 16'haaaa;
            14'h1f88: oData <= 16'hfeaa;
            14'h1f89: oData <= 16'habeb;
            14'h1f8a: oData <= 16'h2bfe;
            14'h1f8b: oData <= 16'h0000;
            14'h1f8c: oData <= 16'h0000;
            14'h1f8d: oData <= 16'h0000;
            14'h1f8e: oData <= 16'h0000;
            14'h1f8f: oData <= 16'h0000;
            14'h1f90: oData <= 16'h0000;
            14'h1f91: oData <= 16'h0000;
            14'h1f92: oData <= 16'h0000;
            14'h1f93: oData <= 16'h0000;
            14'h1f94: oData <= 16'hfea0;
            14'h1f95: oData <= 16'hffff;
            14'h1f96: oData <= 16'hbfeb;
            14'h1f97: oData <= 16'haaaa;
            14'h1f98: oData <= 16'heafa;
            14'h1f99: oData <= 16'hffff;
            14'h1f9a: oData <= 16'hffeb;
            14'h1f9b: oData <= 16'hffaf;
            14'h1f9c: oData <= 16'hfabf;
            14'h1f9d: oData <= 16'habeb;
            14'h1f9e: oData <= 16'h2bfe;
            14'h1f9f: oData <= 16'h0000;
            14'h1fa0: oData <= 16'h0000;
            14'h1fa1: oData <= 16'h0000;
            14'h1fa2: oData <= 16'h0000;
            14'h1fa3: oData <= 16'h0000;
            14'h1fa4: oData <= 16'h0000;
            14'h1fa5: oData <= 16'h0000;
            14'h1fa6: oData <= 16'h0000;
            14'h1fa7: oData <= 16'h0000;
            14'h1fa8: oData <= 16'hfa80;
            14'h1fa9: oData <= 16'hffff;
            14'h1faa: oData <= 16'hbfab;
            14'h1fab: oData <= 16'haabe;
            14'h1fac: oData <= 16'hfaaa;
            14'h1fad: oData <= 16'hffff;
            14'h1fae: oData <= 16'hffeb;
            14'h1faf: oData <= 16'hffaf;
            14'h1fb0: oData <= 16'hfaff;
            14'h1fb1: oData <= 16'haaeb;
            14'h1fb2: oData <= 16'h2bfe;
            14'h1fb3: oData <= 16'h0000;
            14'h1fb4: oData <= 16'h0000;
            14'h1fb5: oData <= 16'h0000;
            14'h1fb6: oData <= 16'h0000;
            14'h1fb7: oData <= 16'h0000;
            14'h1fb8: oData <= 16'h0000;
            14'h1fb9: oData <= 16'h0000;
            14'h1fba: oData <= 16'h0000;
            14'h1fbb: oData <= 16'h0000;
            14'h1fbc: oData <= 16'hea00;
            14'h1fbd: oData <= 16'hffff;
            14'h1fbe: oData <= 16'hbeaf;
            14'h1fbf: oData <= 16'habfe;
            14'h1fc0: oData <= 16'haaaa;
            14'h1fc1: oData <= 16'hffff;
            14'h1fc2: oData <= 16'hffeb;
            14'h1fc3: oData <= 16'hffaf;
            14'h1fc4: oData <= 16'hfaff;
            14'h1fc5: oData <= 16'haaab;
            14'h1fc6: oData <= 16'h2bfe;
            14'h1fc7: oData <= 16'h0000;
            14'h1fc8: oData <= 16'h0000;
            14'h1fc9: oData <= 16'h0000;
            14'h1fca: oData <= 16'h0000;
            14'h1fcb: oData <= 16'h0000;
            14'h1fcc: oData <= 16'h0000;
            14'h1fcd: oData <= 16'h0000;
            14'h1fce: oData <= 16'h0000;
            14'h1fcf: oData <= 16'h0000;
            14'h1fd0: oData <= 16'he800;
            14'h1fd1: oData <= 16'hffff;
            14'h1fd2: oData <= 16'hbabf;
            14'h1fd3: oData <= 16'hbffe;
            14'h1fd4: oData <= 16'haaaa;
            14'h1fd5: oData <= 16'hffaa;
            14'h1fd6: oData <= 16'hffeb;
            14'h1fd7: oData <= 16'hffaf;
            14'h1fd8: oData <= 16'haaab;
            14'h1fd9: oData <= 16'haaaa;
            14'h1fda: oData <= 16'h2bfe;
            14'h1fdb: oData <= 16'h0000;
            14'h1fdc: oData <= 16'h0000;
            14'h1fdd: oData <= 16'h0000;
            14'h1fde: oData <= 16'h0000;
            14'h1fdf: oData <= 16'h0000;
            14'h1fe0: oData <= 16'h0000;
            14'h1fe1: oData <= 16'h0000;
            14'h1fe2: oData <= 16'h0000;
            14'h1fe3: oData <= 16'h0000;
            14'h1fe4: oData <= 16'he800;
            14'h1fe5: oData <= 16'hffff;
            14'h1fe6: oData <= 16'haaff;
            14'h1fe7: oData <= 16'hfffe;
            14'h1fe8: oData <= 16'haabf;
            14'h1fe9: oData <= 16'haaaa;
            14'h1fea: oData <= 16'haaaa;
            14'h1feb: oData <= 16'haaaa;
            14'h1fec: oData <= 16'haaaa;
            14'h1fed: oData <= 16'haaaa;
            14'h1fee: oData <= 16'h2bfe;
            14'h1fef: oData <= 16'h0000;
            14'h1ff0: oData <= 16'h0000;
            14'h1ff1: oData <= 16'h0000;
            14'h1ff2: oData <= 16'h0000;
            14'h1ff3: oData <= 16'h0000;
            14'h1ff4: oData <= 16'h0000;
            14'h1ff5: oData <= 16'h0000;
            14'h1ff6: oData <= 16'h0000;
            14'h1ff7: oData <= 16'h0000;
            14'h1ff8: oData <= 16'ha800;
            14'h1ff9: oData <= 16'hffff;
            14'h1ffa: oData <= 16'habff;
            14'h1ffb: oData <= 16'hffff;
            14'h1ffc: oData <= 16'haebf;
            14'h1ffd: oData <= 16'haaaa;
            14'h1ffe: oData <= 16'haaaa;
            14'h1fff: oData <= 16'haaaa;
            14'h2000: oData <= 16'haaaa;
            14'h2001: oData <= 16'haaaa;
            14'h2002: oData <= 16'h2bfe;
            14'h2003: oData <= 16'h0000;
            14'h2004: oData <= 16'h0000;
            14'h2005: oData <= 16'h0000;
            14'h2006: oData <= 16'h0000;
            14'h2007: oData <= 16'h0000;
            14'h2008: oData <= 16'h0000;
            14'h2009: oData <= 16'h0000;
            14'h200a: oData <= 16'h0000;
            14'h200b: oData <= 16'h0000;
            14'h200c: oData <= 16'ha000;
            14'h200d: oData <= 16'hffff;
            14'h200e: oData <= 16'hafff;
            14'h200f: oData <= 16'hfffe;
            14'h2010: oData <= 16'hfebf;
            14'h2011: oData <= 16'haaab;
            14'h2012: oData <= 16'haaaa;
            14'h2013: oData <= 16'haaaa;
            14'h2014: oData <= 16'haaaa;
            14'h2015: oData <= 16'haaaa;
            14'h2016: oData <= 16'h2bfe;
            14'h2017: oData <= 16'h0000;
            14'h2018: oData <= 16'h0000;
            14'h2019: oData <= 16'h0000;
            14'h201a: oData <= 16'h0000;
            14'h201b: oData <= 16'h0000;
            14'h201c: oData <= 16'h0000;
            14'h201d: oData <= 16'h0000;
            14'h201e: oData <= 16'h0000;
            14'h201f: oData <= 16'h0000;
            14'h2020: oData <= 16'ha000;
            14'h2021: oData <= 16'hfffe;
            14'h2022: oData <= 16'hbfff;
            14'h2023: oData <= 16'hfffa;
            14'h2024: oData <= 16'hfebf;
            14'h2025: oData <= 16'haaff;
            14'h2026: oData <= 16'haaaa;
            14'h2027: oData <= 16'haaaa;
            14'h2028: oData <= 16'haaaa;
            14'h2029: oData <= 16'haaaa;
            14'h202a: oData <= 16'h2bff;
            14'h202b: oData <= 16'h0000;
            14'h202c: oData <= 16'h0000;
            14'h202d: oData <= 16'h0000;
            14'h202e: oData <= 16'h0000;
            14'h202f: oData <= 16'h0000;
            14'h2030: oData <= 16'h0000;
            14'h2031: oData <= 16'h0000;
            14'h2032: oData <= 16'h0000;
            14'h2033: oData <= 16'h0000;
            14'h2034: oData <= 16'h8000;
            14'h2035: oData <= 16'hfffa;
            14'h2036: oData <= 16'hffff;
            14'h2037: oData <= 16'hffaa;
            14'h2038: oData <= 16'hfeaf;
            14'h2039: oData <= 16'hbfff;
            14'h203a: oData <= 16'haaaa;
            14'h203b: oData <= 16'haaaa;
            14'h203c: oData <= 16'haaaa;
            14'h203d: oData <= 16'haeaa;
            14'h203e: oData <= 16'h2bff;
            14'h203f: oData <= 16'h0000;
            14'h2040: oData <= 16'h0000;
            14'h2041: oData <= 16'h0000;
            14'h2042: oData <= 16'h0000;
            14'h2043: oData <= 16'h0000;
            14'h2044: oData <= 16'h0000;
            14'h2045: oData <= 16'h0000;
            14'h2046: oData <= 16'h0000;
            14'h2047: oData <= 16'h0000;
            14'h2048: oData <= 16'h0000;
            14'h2049: oData <= 16'hffea;
            14'h204a: oData <= 16'hffff;
            14'h204b: oData <= 16'hfeab;
            14'h204c: oData <= 16'hffaf;
            14'h204d: oData <= 16'hbfff;
            14'h204e: oData <= 16'haafe;
            14'h204f: oData <= 16'haaaa;
            14'h2050: oData <= 16'haaaa;
            14'h2051: oData <= 16'haebe;
            14'h2052: oData <= 16'h2bff;
            14'h2053: oData <= 16'h0000;
            14'h2054: oData <= 16'h0000;
            14'h2055: oData <= 16'h0000;
            14'h2056: oData <= 16'h0000;
            14'h2057: oData <= 16'h0000;
            14'h2058: oData <= 16'h0000;
            14'h2059: oData <= 16'h0000;
            14'h205a: oData <= 16'h0000;
            14'h205b: oData <= 16'h0000;
            14'h205c: oData <= 16'h0000;
            14'h205d: oData <= 16'hffa8;
            14'h205e: oData <= 16'hffff;
            14'h205f: oData <= 16'heabf;
            14'h2060: oData <= 16'hffaf;
            14'h2061: oData <= 16'hbfff;
            14'h2062: oData <= 16'hfffe;
            14'h2063: oData <= 16'hffab;
            14'h2064: oData <= 16'hafeb;
            14'h2065: oData <= 16'hebaf;
            14'h2066: oData <= 16'h2bff;
            14'h2067: oData <= 16'h0000;
            14'h2068: oData <= 16'h0000;
            14'h2069: oData <= 16'h0000;
            14'h206a: oData <= 16'h0000;
            14'h206b: oData <= 16'h0000;
            14'h206c: oData <= 16'h0000;
            14'h206d: oData <= 16'h0000;
            14'h206e: oData <= 16'h0000;
            14'h206f: oData <= 16'h0000;
            14'h2070: oData <= 16'h0000;
            14'h2071: oData <= 16'hfea8;
            14'h2072: oData <= 16'hffff;
            14'h2073: oData <= 16'haaff;
            14'h2074: oData <= 16'hffaa;
            14'h2075: oData <= 16'hbfff;
            14'h2076: oData <= 16'hfffe;
            14'h2077: oData <= 16'hffeb;
            14'h2078: oData <= 16'habea;
            14'h2079: oData <= 16'heaab;
            14'h207a: oData <= 16'h2bff;
            14'h207b: oData <= 16'h0000;
            14'h207c: oData <= 16'h0000;
            14'h207d: oData <= 16'h0000;
            14'h207e: oData <= 16'h0000;
            14'h207f: oData <= 16'h0000;
            14'h2080: oData <= 16'h0000;
            14'h2081: oData <= 16'h0000;
            14'h2082: oData <= 16'h0000;
            14'h2083: oData <= 16'h0000;
            14'h2084: oData <= 16'h0000;
            14'h2085: oData <= 16'hfa80;
            14'h2086: oData <= 16'hebfe;
            14'h2087: oData <= 16'hafff;
            14'h2088: oData <= 16'hffea;
            14'h2089: oData <= 16'hbfff;
            14'h208a: oData <= 16'hfffe;
            14'h208b: oData <= 16'hffeb;
            14'h208c: oData <= 16'hebfa;
            14'h208d: oData <= 16'hfaef;
            14'h208e: oData <= 16'h2bff;
            14'h208f: oData <= 16'h0000;
            14'h2090: oData <= 16'h0000;
            14'h2091: oData <= 16'h0000;
            14'h2092: oData <= 16'h0000;
            14'h2093: oData <= 16'h0000;
            14'h2094: oData <= 16'h0000;
            14'h2095: oData <= 16'h0000;
            14'h2096: oData <= 16'h0000;
            14'h2097: oData <= 16'h0000;
            14'h2098: oData <= 16'h0000;
            14'h2099: oData <= 16'hea00;
            14'h209a: oData <= 16'hffeb;
            14'h209b: oData <= 16'hfffe;
            14'h209c: oData <= 16'hfaaa;
            14'h209d: oData <= 16'hbfff;
            14'h209e: oData <= 16'hfffe;
            14'h209f: oData <= 16'hbfeb;
            14'h20a0: oData <= 16'heafa;
            14'h20a1: oData <= 16'hfabf;
            14'h20a2: oData <= 16'h2bff;
            14'h20a3: oData <= 16'h0000;
            14'h20a4: oData <= 16'h0000;
            14'h20a5: oData <= 16'h0000;
            14'h20a6: oData <= 16'h0000;
            14'h20a7: oData <= 16'h0000;
            14'h20a8: oData <= 16'h0000;
            14'h20a9: oData <= 16'h0000;
            14'h20aa: oData <= 16'h0000;
            14'h20ab: oData <= 16'h0000;
            14'h20ac: oData <= 16'h0000;
            14'h20ad: oData <= 16'ha800;
            14'h20ae: oData <= 16'hfebf;
            14'h20af: oData <= 16'hffeb;
            14'h20b0: oData <= 16'haaaf;
            14'h20b1: oData <= 16'hbffe;
            14'h20b2: oData <= 16'hfffe;
            14'h20b3: oData <= 16'hbfea;
            14'h20b4: oData <= 16'habfe;
            14'h20b5: oData <= 16'hffaa;
            14'h20b6: oData <= 16'h2bff;
            14'h20b7: oData <= 16'h0000;
            14'h20b8: oData <= 16'h0000;
            14'h20b9: oData <= 16'h0000;
            14'h20ba: oData <= 16'h0000;
            14'h20bb: oData <= 16'h0000;
            14'h20bc: oData <= 16'h0000;
            14'h20bd: oData <= 16'h0000;
            14'h20be: oData <= 16'h0000;
            14'h20bf: oData <= 16'h0000;
            14'h20c0: oData <= 16'h0000;
            14'h20c1: oData <= 16'ha000;
            14'h20c2: oData <= 16'hebfa;
            14'h20c3: oData <= 16'hfebf;
            14'h20c4: oData <= 16'habff;
            14'h20c5: oData <= 16'haaaa;
            14'h20c6: oData <= 16'hfffa;
            14'h20c7: oData <= 16'haffa;
            14'h20c8: oData <= 16'haaaa;
            14'h20c9: oData <= 16'hffea;
            14'h20ca: oData <= 16'habff;
            14'h20cb: oData <= 16'h0000;
            14'h20cc: oData <= 16'h0000;
            14'h20cd: oData <= 16'h0000;
            14'h20ce: oData <= 16'h0000;
            14'h20cf: oData <= 16'h0000;
            14'h20d0: oData <= 16'h0000;
            14'h20d1: oData <= 16'h0000;
            14'h20d2: oData <= 16'h0000;
            14'h20d3: oData <= 16'h0000;
            14'h20d4: oData <= 16'h0000;
            14'h20d5: oData <= 16'h8000;
            14'h20d6: oData <= 16'hbfea;
            14'h20d7: oData <= 16'hebfe;
            14'h20d8: oData <= 16'hffff;
            14'h20d9: oData <= 16'haaaa;
            14'h20da: oData <= 16'haaaa;
            14'h20db: oData <= 16'haaaa;
            14'h20dc: oData <= 16'heaaa;
            14'h20dd: oData <= 16'hffff;
            14'h20de: oData <= 16'habff;
            14'h20df: oData <= 16'h0002;
            14'h20e0: oData <= 16'h0000;
            14'h20e1: oData <= 16'h0000;
            14'h20e2: oData <= 16'h0000;
            14'h20e3: oData <= 16'h0000;
            14'h20e4: oData <= 16'h0000;
            14'h20e5: oData <= 16'h0000;
            14'h20e6: oData <= 16'h0000;
            14'h20e7: oData <= 16'h0000;
            14'h20e8: oData <= 16'h0000;
            14'h20e9: oData <= 16'h0000;
            14'h20ea: oData <= 16'hfea8;
            14'h20eb: oData <= 16'hbfeb;
            14'h20ec: oData <= 16'hfffe;
            14'h20ed: oData <= 16'hffff;
            14'h20ee: oData <= 16'haaab;
            14'h20ef: oData <= 16'heaaa;
            14'h20f0: oData <= 16'hffff;
            14'h20f1: oData <= 16'hffff;
            14'h20f2: oData <= 16'habff;
            14'h20f3: oData <= 16'h0002;
            14'h20f4: oData <= 16'h0000;
            14'h20f5: oData <= 16'h0000;
            14'h20f6: oData <= 16'h0000;
            14'h20f7: oData <= 16'h0000;
            14'h20f8: oData <= 16'h0000;
            14'h20f9: oData <= 16'h0000;
            14'h20fa: oData <= 16'h0000;
            14'h20fb: oData <= 16'h0000;
            14'h20fc: oData <= 16'h0000;
            14'h20fd: oData <= 16'h0000;
            14'h20fe: oData <= 16'heaa0;
            14'h20ff: oData <= 16'hfebf;
            14'h2100: oData <= 16'hffab;
            14'h2101: oData <= 16'hffff;
            14'h2102: oData <= 16'hffff;
            14'h2103: oData <= 16'hffff;
            14'h2104: oData <= 16'hffff;
            14'h2105: oData <= 16'hfeff;
            14'h2106: oData <= 16'habff;
            14'h2107: oData <= 16'h0002;
            14'h2108: oData <= 16'h0000;
            14'h2109: oData <= 16'h0000;
            14'h210a: oData <= 16'h0000;
            14'h210b: oData <= 16'h0000;
            14'h210c: oData <= 16'h0000;
            14'h210d: oData <= 16'h0000;
            14'h210e: oData <= 16'h0000;
            14'h210f: oData <= 16'h0000;
            14'h2110: oData <= 16'h0000;
            14'h2111: oData <= 16'h0000;
            14'h2112: oData <= 16'haa00;
            14'h2113: oData <= 16'hebfe;
            14'h2114: oData <= 16'heaff;
            14'h2115: oData <= 16'hffff;
            14'h2116: oData <= 16'hffff;
            14'h2117: oData <= 16'hffff;
            14'h2118: oData <= 16'hffff;
            14'h2119: oData <= 16'hffbf;
            14'h211a: oData <= 16'haffe;
            14'h211b: oData <= 16'h0000;
            14'h211c: oData <= 16'h0000;
            14'h211d: oData <= 16'h0000;
            14'h211e: oData <= 16'h0000;
            14'h211f: oData <= 16'h0000;
            14'h2120: oData <= 16'h0000;
            14'h2121: oData <= 16'h0000;
            14'h2122: oData <= 16'h0000;
            14'h2123: oData <= 16'h0000;
            14'h2124: oData <= 16'h0000;
            14'h2125: oData <= 16'h0000;
            14'h2126: oData <= 16'ha000;
            14'h2127: oData <= 16'hbfea;
            14'h2128: oData <= 16'hbffa;
            14'h2129: oData <= 16'hfffe;
            14'h212a: oData <= 16'haaab;
            14'h212b: oData <= 16'haaaa;
            14'h212c: oData <= 16'hfffe;
            14'h212d: oData <= 16'hffeb;
            14'h212e: oData <= 16'haffe;
            14'h212f: oData <= 16'h0000;
            14'h2130: oData <= 16'h0000;
            14'h2131: oData <= 16'h0000;
            14'h2132: oData <= 16'h0000;
            14'h2133: oData <= 16'h0000;
            14'h2134: oData <= 16'h0000;
            14'h2135: oData <= 16'h0000;
            14'h2136: oData <= 16'h0000;
            14'h2137: oData <= 16'h0000;
            14'h2138: oData <= 16'h0000;
            14'h2139: oData <= 16'h0000;
            14'h213a: oData <= 16'h0000;
            14'h213b: oData <= 16'hfeaa;
            14'h213c: oData <= 16'hfeaf;
            14'h213d: oData <= 16'hfaab;
            14'h213e: oData <= 16'hffff;
            14'h213f: oData <= 16'hffff;
            14'h2140: oData <= 16'hffff;
            14'h2141: oData <= 16'hfffe;
            14'h2142: oData <= 16'haffe;
            14'h2143: oData <= 16'h0000;
            14'h2144: oData <= 16'h0000;
            14'h2145: oData <= 16'h0000;
            14'h2146: oData <= 16'h0000;
            14'h2147: oData <= 16'h0000;
            14'h2148: oData <= 16'h0000;
            14'h2149: oData <= 16'h0a00;
            14'h214a: oData <= 16'h0000;
            14'h214b: oData <= 16'h0000;
            14'h214c: oData <= 16'h0000;
            14'h214d: oData <= 16'h0000;
            14'h214e: oData <= 16'h0000;
            14'h214f: oData <= 16'haaa0;
            14'h2150: oData <= 16'habff;
            14'h2151: oData <= 16'hafff;
            14'h2152: oData <= 16'haaaa;
            14'h2153: oData <= 16'hfffe;
            14'h2154: oData <= 16'haaff;
            14'h2155: oData <= 16'hbfff;
            14'h2156: oData <= 16'hafff;
            14'h2157: oData <= 16'h0000;
            14'h2158: oData <= 16'h0000;
            14'h2159: oData <= 16'h0000;
            14'h215a: oData <= 16'h0000;
            14'h215b: oData <= 16'h0000;
            14'h215c: oData <= 16'h0000;
            14'h215d: oData <= 16'h2a80;
            14'h215e: oData <= 16'h0000;
            14'h215f: oData <= 16'h0000;
            14'h2160: oData <= 16'h0000;
            14'h2161: oData <= 16'h0000;
            14'h2162: oData <= 16'h0000;
            14'h2163: oData <= 16'haa00;
            14'h2164: oData <= 16'hfffa;
            14'h2165: oData <= 16'hfeaa;
            14'h2166: oData <= 16'hffff;
            14'h2167: oData <= 16'haaab;
            14'h2168: oData <= 16'hffaa;
            14'h2169: oData <= 16'hebff;
            14'h216a: oData <= 16'hafff;
            14'h216b: oData <= 16'h0000;
            14'h216c: oData <= 16'h0000;
            14'h216d: oData <= 16'h0000;
            14'h216e: oData <= 16'h0000;
            14'h216f: oData <= 16'h0000;
            14'h2170: oData <= 16'h0000;
            14'h2171: oData <= 16'h2aa0;
            14'h2172: oData <= 16'h0000;
            14'h2173: oData <= 16'h0000;
            14'h2174: oData <= 16'h0000;
            14'h2175: oData <= 16'h0000;
            14'h2176: oData <= 16'h0000;
            14'h2177: oData <= 16'h8000;
            14'h2178: oData <= 16'hffaa;
            14'h2179: oData <= 16'habff;
            14'h217a: oData <= 16'hffea;
            14'h217b: oData <= 16'hffff;
            14'h217c: oData <= 16'hffff;
            14'h217d: oData <= 16'hfeff;
            14'h217e: oData <= 16'hafff;
            14'h217f: oData <= 16'h0000;
            14'h2180: oData <= 16'h0000;
            14'h2181: oData <= 16'h0000;
            14'h2182: oData <= 16'h0000;
            14'h2183: oData <= 16'h0000;
            14'h2184: oData <= 16'h0000;
            14'h2185: oData <= 16'h2aa0;
            14'h2186: oData <= 16'h0000;
            14'h2187: oData <= 16'h0000;
            14'h2188: oData <= 16'h0000;
            14'h2189: oData <= 16'h0000;
            14'h218a: oData <= 16'h0000;
            14'h218b: oData <= 16'h0000;
            14'h218c: oData <= 16'hfaa8;
            14'h218d: oData <= 16'hffff;
            14'h218e: oData <= 16'haabf;
            14'h218f: oData <= 16'hfeaa;
            14'h2190: oData <= 16'hffff;
            14'h2191: oData <= 16'hffaa;
            14'h2192: oData <= 16'habff;
            14'h2193: oData <= 16'h0000;
            14'h2194: oData <= 16'h0000;
            14'h2195: oData <= 16'h0000;
            14'h2196: oData <= 16'h0000;
            14'h2197: oData <= 16'h0000;
            14'h2198: oData <= 16'h0000;
            14'h2199: oData <= 16'h0aa8;
            14'h219a: oData <= 16'h0000;
            14'h219b: oData <= 16'h0000;
            14'h219c: oData <= 16'h0000;
            14'h219d: oData <= 16'h0000;
            14'h219e: oData <= 16'h0000;
            14'h219f: oData <= 16'h0000;
            14'h21a0: oData <= 16'haa80;
            14'h21a1: oData <= 16'hffff;
            14'h21a2: oData <= 16'hffff;
            14'h21a3: oData <= 16'habff;
            14'h21a4: oData <= 16'haaaa;
            14'h21a5: oData <= 16'hffff;
            14'h21a6: oData <= 16'h2bff;
            14'h21a7: oData <= 16'h0000;
            14'h21a8: oData <= 16'h0000;
            14'h21a9: oData <= 16'h0000;
            14'h21aa: oData <= 16'h0000;
            14'h21ab: oData <= 16'h0000;
            14'h21ac: oData <= 16'h0000;
            14'h21ad: oData <= 16'h0aa8;
            14'h21ae: oData <= 16'h0000;
            14'h21af: oData <= 16'h0000;
            14'h21b0: oData <= 16'h0000;
            14'h21b1: oData <= 16'h0000;
            14'h21b2: oData <= 16'h0000;
            14'h21b3: oData <= 16'h0000;
            14'h21b4: oData <= 16'ha800;
            14'h21b5: oData <= 16'hfffa;
            14'h21b6: oData <= 16'hffff;
            14'h21b7: oData <= 16'hffff;
            14'h21b8: oData <= 16'hffff;
            14'h21b9: oData <= 16'hffff;
            14'h21ba: oData <= 16'h2aff;
            14'h21bb: oData <= 16'h0000;
            14'h21bc: oData <= 16'h0000;
            14'h21bd: oData <= 16'h0000;
            14'h21be: oData <= 16'h0000;
            14'h21bf: oData <= 16'h0000;
            14'h21c0: oData <= 16'h0000;
            14'h21c1: oData <= 16'h02aa;
            14'h21c2: oData <= 16'h0000;
            14'h21c3: oData <= 16'h0000;
            14'h21c4: oData <= 16'h0000;
            14'h21c5: oData <= 16'h0000;
            14'h21c6: oData <= 16'h0000;
            14'h21c7: oData <= 16'h0000;
            14'h21c8: oData <= 16'h8000;
            14'h21c9: oData <= 16'hffaa;
            14'h21ca: oData <= 16'hffff;
            14'h21cb: oData <= 16'hffff;
            14'h21cc: oData <= 16'hffff;
            14'h21cd: oData <= 16'hffff;
            14'h21ce: oData <= 16'h0aff;
            14'h21cf: oData <= 16'h0000;
            14'h21d0: oData <= 16'h0000;
            14'h21d1: oData <= 16'h0000;
            14'h21d2: oData <= 16'h0000;
            14'h21d3: oData <= 16'h0000;
            14'h21d4: oData <= 16'h0000;
            14'h21d5: oData <= 16'h02aa;
            14'h21d6: oData <= 16'h0000;
            14'h21d7: oData <= 16'h0000;
            14'h21d8: oData <= 16'h0000;
            14'h21d9: oData <= 16'h0000;
            14'h21da: oData <= 16'h0000;
            14'h21db: oData <= 16'h0000;
            14'h21dc: oData <= 16'h0000;
            14'h21dd: oData <= 16'haaa8;
            14'h21de: oData <= 16'hfffe;
            14'h21df: oData <= 16'hffff;
            14'h21e0: oData <= 16'hffff;
            14'h21e1: oData <= 16'hffff;
            14'h21e2: oData <= 16'h0abf;
            14'h21e3: oData <= 16'h0000;
            14'h21e4: oData <= 16'h0000;
            14'h21e5: oData <= 16'h0000;
            14'h21e6: oData <= 16'h0000;
            14'h21e7: oData <= 16'h0000;
            14'h21e8: oData <= 16'h0000;
            14'h21e9: oData <= 16'h00aa;
            14'h21ea: oData <= 16'h0000;
            14'h21eb: oData <= 16'h02a8;
            14'h21ec: oData <= 16'h0000;
            14'h21ed: oData <= 16'h0000;
            14'h21ee: oData <= 16'h0000;
            14'h21ef: oData <= 16'h0000;
            14'h21f0: oData <= 16'h0000;
            14'h21f1: oData <= 16'haa80;
            14'h21f2: oData <= 16'hfeaa;
            14'h21f3: oData <= 16'hffff;
            14'h21f4: oData <= 16'hffff;
            14'h21f5: oData <= 16'hffff;
            14'h21f6: oData <= 16'h02ab;
            14'h21f7: oData <= 16'h0000;
            14'h21f8: oData <= 16'h0000;
            14'h21f9: oData <= 16'h0000;
            14'h21fa: oData <= 16'h0000;
            14'h21fb: oData <= 16'h0000;
            14'h21fc: oData <= 16'h8000;
            14'h21fd: oData <= 16'h00aa;
            14'h21fe: oData <= 16'h0000;
            14'h21ff: oData <= 16'h0aaa;
            14'h2200: oData <= 16'h0000;
            14'h2201: oData <= 16'h0000;
            14'h2202: oData <= 16'h0000;
            14'h2203: oData <= 16'h0000;
            14'h2204: oData <= 16'h0000;
            14'h2205: oData <= 16'haa00;
            14'h2206: oData <= 16'haaaa;
            14'h2207: oData <= 16'hfffe;
            14'h2208: oData <= 16'hffff;
            14'h2209: oData <= 16'hffff;
            14'h220a: oData <= 16'h00aa;
            14'h220b: oData <= 16'h0000;
            14'h220c: oData <= 16'h0000;
            14'h220d: oData <= 16'h0000;
            14'h220e: oData <= 16'h0000;
            14'h220f: oData <= 16'h0000;
            14'h2210: oData <= 16'h8000;
            14'h2211: oData <= 16'h00aa;
            14'h2212: oData <= 16'h8000;
            14'h2213: oData <= 16'h0aaa;
            14'h2214: oData <= 16'h0000;
            14'h2215: oData <= 16'h0000;
            14'h2216: oData <= 16'h0000;
            14'h2217: oData <= 16'h0000;
            14'h2218: oData <= 16'h0000;
            14'h2219: oData <= 16'haa00;
            14'h221a: oData <= 16'haa0a;
            14'h221b: oData <= 16'hfeaa;
            14'h221c: oData <= 16'hffff;
            14'h221d: oData <= 16'habff;
            14'h221e: oData <= 16'h000a;
            14'h221f: oData <= 16'h0000;
            14'h2220: oData <= 16'h0000;
            14'h2221: oData <= 16'h0000;
            14'h2222: oData <= 16'h0000;
            14'h2223: oData <= 16'h0000;
            14'h2224: oData <= 16'h8000;
            14'h2225: oData <= 16'h002a;
            14'h2226: oData <= 16'ha000;
            14'h2227: oData <= 16'h2aaa;
            14'h2228: oData <= 16'h0000;
            14'h2229: oData <= 16'h0000;
            14'h222a: oData <= 16'h0000;
            14'h222b: oData <= 16'h0000;
            14'h222c: oData <= 16'h0000;
            14'h222d: oData <= 16'ha800;
            14'h222e: oData <= 16'h000a;
            14'h222f: oData <= 16'haaaa;
            14'h2230: oData <= 16'haaaa;
            14'h2231: oData <= 16'haaaa;
            14'h2232: oData <= 16'h0000;
            14'h2233: oData <= 16'h0000;
            14'h2234: oData <= 16'h0000;
            14'h2235: oData <= 16'h0000;
            14'h2236: oData <= 16'h0000;
            14'h2237: oData <= 16'h0000;
            14'h2238: oData <= 16'ha000;
            14'h2239: oData <= 16'h002a;
            14'h223a: oData <= 16'ha800;
            14'h223b: oData <= 16'h2aaa;
            14'h223c: oData <= 16'h0000;
            14'h223d: oData <= 16'h0000;
            14'h223e: oData <= 16'h0000;
            14'h223f: oData <= 16'h0000;
            14'h2240: oData <= 16'h0000;
            14'h2241: oData <= 16'ha800;
            14'h2242: oData <= 16'h000a;
            14'h2243: oData <= 16'haa00;
            14'h2244: oData <= 16'haaaa;
            14'h2245: oData <= 16'h0aaa;
            14'h2246: oData <= 16'h02a0;
            14'h2247: oData <= 16'h0000;
            14'h2248: oData <= 16'h0000;
            14'h2249: oData <= 16'h0000;
            14'h224a: oData <= 16'h0000;
            14'h224b: oData <= 16'h0000;
            14'h224c: oData <= 16'ha000;
            14'h224d: oData <= 16'h002a;
            14'h224e: oData <= 16'ha800;
            14'h224f: oData <= 16'h2a8a;
            14'h2250: oData <= 16'h2800;
            14'h2251: oData <= 16'h0000;
            14'h2252: oData <= 16'h0000;
            14'h2253: oData <= 16'h0000;
            14'h2254: oData <= 16'h0000;
            14'h2255: oData <= 16'ha800;
            14'h2256: oData <= 16'h000a;
            14'h2257: oData <= 16'h8000;
            14'h2258: oData <= 16'haaaa;
            14'h2259: oData <= 16'h0aaa;
            14'h225a: oData <= 16'h0aa8;
            14'h225b: oData <= 16'h0000;
            14'h225c: oData <= 16'h0000;
            14'h225d: oData <= 16'h0000;
            14'h225e: oData <= 16'h0000;
            14'h225f: oData <= 16'h0000;
            14'h2260: oData <= 16'ha000;
            14'h2261: oData <= 16'h000a;
            14'h2262: oData <= 16'ha800;
            14'h2263: oData <= 16'h2a82;
            14'h2264: oData <= 16'haa00;
            14'h2265: oData <= 16'h0000;
            14'h2266: oData <= 16'h0000;
            14'h2267: oData <= 16'h0000;
            14'h2268: oData <= 16'h0000;
            14'h2269: oData <= 16'ha800;
            14'h226a: oData <= 16'h002a;
            14'h226b: oData <= 16'haa00;
            14'h226c: oData <= 16'haaaa;
            14'h226d: oData <= 16'h02aa;
            14'h226e: oData <= 16'h0aa8;
            14'h226f: oData <= 16'h0000;
            14'h2270: oData <= 16'h0000;
            14'h2271: oData <= 16'h0000;
            14'h2272: oData <= 16'h0000;
            14'h2273: oData <= 16'h0000;
            14'h2274: oData <= 16'ha000;
            14'h2275: oData <= 16'h000a;
            14'h2276: oData <= 16'haa00;
            14'h2277: oData <= 16'h2a82;
            14'h2278: oData <= 16'haa80;
            14'h2279: oData <= 16'h0000;
            14'h227a: oData <= 16'h0000;
            14'h227b: oData <= 16'h0000;
            14'h227c: oData <= 16'h0000;
            14'h227d: oData <= 16'ha000;
            14'h227e: oData <= 16'h002a;
            14'h227f: oData <= 16'haaaa;
            14'h2280: oData <= 16'haaaa;
            14'h2281: oData <= 16'h00aa;
            14'h2282: oData <= 16'h0aaa;
            14'h2283: oData <= 16'h0000;
            14'h2284: oData <= 16'h0000;
            14'h2285: oData <= 16'h0000;
            14'h2286: oData <= 16'h0000;
            14'h2287: oData <= 16'h0000;
            14'h2288: oData <= 16'ha000;
            14'h2289: oData <= 16'h002a;
            14'h228a: oData <= 16'haa00;
            14'h228b: oData <= 16'h2a82;
            14'h228c: oData <= 16'haa80;
            14'h228d: oData <= 16'h0000;
            14'h228e: oData <= 16'h0000;
            14'h228f: oData <= 16'h0000;
            14'h2290: oData <= 16'h0000;
            14'h2291: oData <= 16'ha000;
            14'h2292: oData <= 16'haa2a;
            14'h2293: oData <= 16'haaaa;
            14'h2294: oData <= 16'haaaa;
            14'h2295: oData <= 16'h0000;
            14'h2296: oData <= 16'h02aa;
            14'h2297: oData <= 16'h0000;
            14'h2298: oData <= 16'h0000;
            14'h2299: oData <= 16'h0000;
            14'h229a: oData <= 16'h0000;
            14'h229b: oData <= 16'h0000;
            14'h229c: oData <= 16'ha000;
            14'h229d: oData <= 16'h00aa;
            14'h229e: oData <= 16'haa00;
            14'h229f: oData <= 16'h2a80;
            14'h22a0: oData <= 16'h2aa0;
            14'h22a1: oData <= 16'h0000;
            14'h22a2: oData <= 16'h0000;
            14'h22a3: oData <= 16'h0000;
            14'h22a4: oData <= 16'h0000;
            14'h22a5: oData <= 16'ha000;
            14'h22a6: oData <= 16'haaaa;
            14'h22a7: oData <= 16'haaaa;
            14'h22a8: oData <= 16'h00aa;
            14'h22a9: oData <= 16'h8000;
            14'h22aa: oData <= 16'h02aa;
            14'h22ab: oData <= 16'h0000;
            14'h22ac: oData <= 16'h0000;
            14'h22ad: oData <= 16'h0000;
            14'h22ae: oData <= 16'h0000;
            14'h22af: oData <= 16'h0000;
            14'h22b0: oData <= 16'ha000;
            14'h22b1: oData <= 16'h02aa;
            14'h22b2: oData <= 16'haa00;
            14'h22b3: oData <= 16'h2a80;
            14'h22b4: oData <= 16'h2aa0;
            14'h22b5: oData <= 16'h0000;
            14'h22b6: oData <= 16'h0000;
            14'h22b7: oData <= 16'h0000;
            14'h22b8: oData <= 16'h0000;
            14'h22b9: oData <= 16'ha000;
            14'h22ba: oData <= 16'haaaa;
            14'h22bb: oData <= 16'haaaa;
            14'h22bc: oData <= 16'h0000;
            14'h22bd: oData <= 16'h8000;
            14'h22be: oData <= 16'h00aa;
            14'h22bf: oData <= 16'h0000;
            14'h22c0: oData <= 16'h0000;
            14'h22c1: oData <= 16'h0000;
            14'h22c2: oData <= 16'h0000;
            14'h22c3: oData <= 16'h0000;
            14'h22c4: oData <= 16'h8000;
            14'h22c5: oData <= 16'h0aaa;
            14'h22c6: oData <= 16'haa80;
            14'h22c7: oData <= 16'h2aa0;
            14'h22c8: oData <= 16'h0aa8;
            14'h22c9: oData <= 16'h0000;
            14'h22ca: oData <= 16'h0000;
            14'h22cb: oData <= 16'h0000;
            14'h22cc: oData <= 16'h0000;
            14'h22cd: oData <= 16'ha800;
            14'h22ce: oData <= 16'haaaa;
            14'h22cf: oData <= 16'h02aa;
            14'h22d0: oData <= 16'h0000;
            14'h22d1: oData <= 16'ha000;
            14'h22d2: oData <= 16'h00aa;
            14'h22d3: oData <= 16'h0000;
            14'h22d4: oData <= 16'h0000;
            14'h22d5: oData <= 16'h0000;
            14'h22d6: oData <= 16'h0000;
            14'h22d7: oData <= 16'h0000;
            14'h22d8: oData <= 16'h0000;
            14'h22d9: oData <= 16'h0aaa;
            14'h22da: oData <= 16'haa80;
            14'h22db: oData <= 16'h2aa0;
            14'h22dc: oData <= 16'h0aa8;
            14'h22dd: oData <= 16'h0000;
            14'h22de: oData <= 16'h0000;
            14'h22df: oData <= 16'h0000;
            14'h22e0: oData <= 16'h0000;
            14'h22e1: oData <= 16'haa80;
            14'h22e2: oData <= 16'haaaa;
            14'h22e3: oData <= 16'h0002;
            14'h22e4: oData <= 16'h0000;
            14'h22e5: oData <= 16'ha000;
            14'h22e6: oData <= 16'h002a;
            14'h22e7: oData <= 16'h0000;
            14'h22e8: oData <= 16'h0000;
            14'h22e9: oData <= 16'h0000;
            14'h22ea: oData <= 16'h0000;
            14'h22eb: oData <= 16'h0000;
            14'h22ec: oData <= 16'h0000;
            14'h22ed: oData <= 16'haaa0;
            14'h22ee: oData <= 16'h2a80;
            14'h22ef: oData <= 16'h0aa8;
            14'h22f0: oData <= 16'h02aa;
            14'h22f1: oData <= 16'h0000;
            14'h22f2: oData <= 16'h0000;
            14'h22f3: oData <= 16'h0000;
            14'h22f4: oData <= 16'h0000;
            14'h22f5: oData <= 16'haaa8;
            14'h22f6: oData <= 16'h02aa;
            14'h22f7: oData <= 16'h0000;
            14'h22f8: oData <= 16'h0000;
            14'h22f9: oData <= 16'ha800;
            14'h22fa: oData <= 16'h002a;
            14'h22fb: oData <= 16'h0000;
            14'h22fc: oData <= 16'h0000;
            14'h22fd: oData <= 16'h0000;
            14'h22fe: oData <= 16'h0000;
            14'h22ff: oData <= 16'h0000;
            14'h2300: oData <= 16'h0000;
            14'h2301: oData <= 16'haaa0;
            14'h2302: oData <= 16'haa82;
            14'h2303: oData <= 16'h0aaa;
            14'h2304: oData <= 16'h02aa;
            14'h2305: oData <= 16'h0000;
            14'h2306: oData <= 16'h0000;
            14'h2307: oData <= 16'h0000;
            14'h2308: oData <= 16'h8000;
            14'h2309: oData <= 16'haaaa;
            14'h230a: oData <= 16'h02aa;
            14'h230b: oData <= 16'h0000;
            14'h230c: oData <= 16'h0000;
            14'h230d: oData <= 16'ha800;
            14'h230e: oData <= 16'h000a;
            14'h230f: oData <= 16'h0000;
            14'h2310: oData <= 16'h0000;
            14'h2311: oData <= 16'h0000;
            14'h2312: oData <= 16'h0000;
            14'h2313: oData <= 16'h0000;
            14'h2314: oData <= 16'h0000;
            14'h2315: oData <= 16'haa80;
            14'h2316: oData <= 16'haa82;
            14'h2317: oData <= 16'h0aaa;
            14'h2318: oData <= 16'h00aa;
            14'h2319: oData <= 16'h0000;
            14'h231a: oData <= 16'h0000;
            14'h231b: oData <= 16'h0000;
            14'h231c: oData <= 16'ha800;
            14'h231d: oData <= 16'haaaa;
            14'h231e: oData <= 16'h02aa;
            14'h231f: oData <= 16'h0000;
            14'h2320: oData <= 16'h0000;
            14'h2321: oData <= 16'ha800;
            14'h2322: oData <= 16'h000a;
            14'h2323: oData <= 16'h0000;
            14'h2324: oData <= 16'h0000;
            14'h2325: oData <= 16'h0000;
            14'h2326: oData <= 16'h0000;
            14'h2327: oData <= 16'h0000;
            14'h2328: oData <= 16'h0000;
            14'h2329: oData <= 16'haa00;
            14'h232a: oData <= 16'haa80;
            14'h232b: oData <= 16'h82aa;
            14'h232c: oData <= 16'h00aa;
            14'h232d: oData <= 16'h0000;
            14'h232e: oData <= 16'h0000;
            14'h232f: oData <= 16'h0000;
            14'h2330: oData <= 16'haa80;
            14'h2331: oData <= 16'h0aaa;
            14'h2332: oData <= 16'h02aa;
            14'h2333: oData <= 16'h0000;
            14'h2334: oData <= 16'h0000;
            14'h2335: oData <= 16'haa00;
            14'h2336: oData <= 16'h000a;
            14'h2337: oData <= 16'h0000;
            14'h2338: oData <= 16'h0000;
            14'h2339: oData <= 16'h0000;
            14'h233a: oData <= 16'h0000;
            14'h233b: oData <= 16'h0000;
            14'h233c: oData <= 16'h0000;
            14'h233d: oData <= 16'h0000;
            14'h233e: oData <= 16'haa00;
            14'h233f: oData <= 16'h802a;
            14'h2340: oData <= 16'h00aa;
            14'h2341: oData <= 16'h0000;
            14'h2342: oData <= 16'h0000;
            14'h2343: oData <= 16'h0000;
            14'h2344: oData <= 16'haaa8;
            14'h2345: oData <= 16'h00aa;
            14'h2346: oData <= 16'h02aa;
            14'h2347: oData <= 16'h0000;
            14'h2348: oData <= 16'h0000;
            14'h2349: oData <= 16'haa00;
            14'h234a: oData <= 16'h0002;
            14'h234b: oData <= 16'h0000;
            14'h234c: oData <= 16'h0000;
            14'h234d: oData <= 16'h0000;
            14'h234e: oData <= 16'h0000;
            14'h234f: oData <= 16'h0000;
            14'h2350: oData <= 16'h0000;
            14'h2351: oData <= 16'h0000;
            14'h2352: oData <= 16'ha000;
            14'h2353: oData <= 16'h8002;
            14'h2354: oData <= 16'h002a;
            14'h2355: oData <= 16'h0000;
            14'h2356: oData <= 16'h0000;
            14'h2357: oData <= 16'ha000;
            14'h2358: oData <= 16'haaaa;
            14'h2359: oData <= 16'h000a;
            14'h235a: oData <= 16'h0aaa;
            14'h235b: oData <= 16'h0000;
            14'h235c: oData <= 16'h0000;
            14'h235d: oData <= 16'haa80;
            14'h235e: oData <= 16'h0002;
            14'h235f: oData <= 16'h0000;
            14'h2360: oData <= 16'h0000;
            14'h2361: oData <= 16'h0000;
            14'h2362: oData <= 16'h0000;
            14'h2363: oData <= 16'h0000;
            14'h2364: oData <= 16'h0000;
            14'h2365: oData <= 16'h0000;
            14'h2366: oData <= 16'h0000;
            14'h2367: oData <= 16'ha000;
            14'h2368: oData <= 16'h002a;
            14'h2369: oData <= 16'h0000;
            14'h236a: oData <= 16'ha000;
            14'h236b: oData <= 16'haaaa;
            14'h236c: oData <= 16'haaaa;
            14'h236d: oData <= 16'h0000;
            14'h236e: oData <= 16'h0aa8;
            14'h236f: oData <= 16'h0000;
            14'h2370: oData <= 16'h0000;
            14'h2371: oData <= 16'haa80;
            14'h2372: oData <= 16'h0000;
            14'h2373: oData <= 16'h0000;
            14'h2374: oData <= 16'h0000;
            14'h2375: oData <= 16'h0000;
            14'h2376: oData <= 16'h0000;
            14'h2377: oData <= 16'h0000;
            14'h2378: oData <= 16'h0000;
            14'h2379: oData <= 16'h0000;
            14'h237a: oData <= 16'h0000;
            14'h237b: oData <= 16'ha000;
            14'h237c: oData <= 16'h002a;
            14'h237d: oData <= 16'ha800;
            14'h237e: oData <= 16'haaaa;
            14'h237f: oData <= 16'haaaa;
            14'h2380: oData <= 16'h0aaa;
            14'h2381: oData <= 16'h0000;
            14'h2382: oData <= 16'h0aa8;
            14'h2383: oData <= 16'h0000;
            14'h2384: oData <= 16'h0000;
            14'h2385: oData <= 16'haaa0;
            14'h2386: oData <= 16'h0000;
            14'h2387: oData <= 16'h0000;
            14'h2388: oData <= 16'h0000;
            14'h2389: oData <= 16'h0000;
            14'h238a: oData <= 16'h0000;
            14'h238b: oData <= 16'h0000;
            14'h238c: oData <= 16'h0000;
            14'h238d: oData <= 16'h0000;
            14'h238e: oData <= 16'h0000;
            14'h238f: oData <= 16'ha000;
            14'h2390: oData <= 16'h000a;
            14'h2391: oData <= 16'haa00;
            14'h2392: oData <= 16'haaaa;
            14'h2393: oData <= 16'haaaa;
            14'h2394: oData <= 16'h00aa;
            14'h2395: oData <= 16'h0000;
            14'h2396: oData <= 16'h0aa8;
            14'h2397: oData <= 16'h0000;
            14'h2398: oData <= 16'h0000;
            14'h2399: oData <= 16'h2aa8;
            14'h239a: oData <= 16'h0000;
            14'h239b: oData <= 16'h0000;
            14'h239c: oData <= 16'h0000;
            14'h239d: oData <= 16'h0000;
            14'h239e: oData <= 16'h0000;
            14'h239f: oData <= 16'h0000;
            14'h23a0: oData <= 16'h0000;
            14'h23a1: oData <= 16'h0000;
            14'h23a2: oData <= 16'h0000;
            14'h23a3: oData <= 16'ha800;
            14'h23a4: oData <= 16'h000a;
            14'h23a5: oData <= 16'haa00;
            14'h23a6: oData <= 16'haaaa;
            14'h23a7: oData <= 16'haaaa;
            14'h23a8: oData <= 16'h000a;
            14'h23a9: oData <= 16'h0000;
            14'h23aa: oData <= 16'h2aa8;
            14'h23ab: oData <= 16'h0000;
            14'h23ac: oData <= 16'ha000;
            14'h23ad: oData <= 16'h2aaa;
            14'h23ae: oData <= 16'h0000;
            14'h23af: oData <= 16'h0000;
            14'h23b0: oData <= 16'h0000;
            14'h23b1: oData <= 16'h0000;
            14'h23b2: oData <= 16'h0000;
            14'h23b3: oData <= 16'h0000;
            14'h23b4: oData <= 16'h0000;
            14'h23b5: oData <= 16'h0000;
            14'h23b6: oData <= 16'h0000;
            14'h23b7: oData <= 16'ha800;
            14'h23b8: oData <= 16'h000a;
            14'h23b9: oData <= 16'haa00;
            14'h23ba: oData <= 16'haaaa;
            14'h23bb: oData <= 16'haaaa;
            14'h23bc: oData <= 16'h0000;
            14'h23bd: oData <= 16'h0000;
            14'h23be: oData <= 16'h2aa0;
            14'h23bf: oData <= 16'h0000;
            14'h23c0: oData <= 16'haa80;
            14'h23c1: oData <= 16'h2aaa;
            14'h23c2: oData <= 16'h0000;
            14'h23c3: oData <= 16'h0000;
            14'h23c4: oData <= 16'h0000;
            14'h23c5: oData <= 16'h0000;
            14'h23c6: oData <= 16'h0000;
            14'h23c7: oData <= 16'h0000;
            14'h23c8: oData <= 16'h0000;
            14'h23c9: oData <= 16'h0000;
            14'h23ca: oData <= 16'h0000;
            14'h23cb: oData <= 16'ha800;
            14'h23cc: oData <= 16'h0002;
            14'h23cd: oData <= 16'ha800;
            14'h23ce: oData <= 16'h2aaa;
            14'h23cf: oData <= 16'h0000;
            14'h23d0: oData <= 16'h0000;
            14'h23d1: oData <= 16'h0000;
            14'h23d2: oData <= 16'h2aa0;
            14'h23d3: oData <= 16'h0000;
            14'h23d4: oData <= 16'haaaa;
            14'h23d5: oData <= 16'h0aaa;
            14'h23d6: oData <= 16'h0000;
            14'h23d7: oData <= 16'h0000;
            14'h23d8: oData <= 16'h0000;
            14'h23d9: oData <= 16'h0000;
            14'h23da: oData <= 16'h0000;
            14'h23db: oData <= 16'h0000;
            14'h23dc: oData <= 16'h0000;
            14'h23dd: oData <= 16'h0000;
            14'h23de: oData <= 16'h0000;
            14'h23df: oData <= 16'ha800;
            14'h23e0: oData <= 16'h000a;
            14'h23e1: oData <= 16'h0000;
            14'h23e2: oData <= 16'h0000;
            14'h23e3: oData <= 16'ha000;
            14'h23e4: oData <= 16'h0002;
            14'h23e5: oData <= 16'h0000;
            14'h23e6: oData <= 16'h2aa0;
            14'h23e7: oData <= 16'ha800;
            14'h23e8: oData <= 16'haaaa;
            14'h23e9: oData <= 16'h02aa;
            14'h23ea: oData <= 16'h0000;
            14'h23eb: oData <= 16'h0000;
            14'h23ec: oData <= 16'h0000;
            14'h23ed: oData <= 16'h0000;
            14'h23ee: oData <= 16'h0000;
            14'h23ef: oData <= 16'h0000;
            14'h23f0: oData <= 16'h0000;
            14'h23f1: oData <= 16'h0000;
            14'h23f2: oData <= 16'h0000;
            14'h23f3: oData <= 16'ha800;
            14'h23f4: oData <= 16'h00aa;
            14'h23f5: oData <= 16'h0000;
            14'h23f6: oData <= 16'h0000;
            14'h23f7: oData <= 16'ha800;
            14'h23f8: oData <= 16'h2aaa;
            14'h23f9: oData <= 16'h0000;
            14'h23fa: oData <= 16'haaa0;
            14'h23fb: oData <= 16'haaa0;
            14'h23fc: oData <= 16'haaaa;
            14'h23fd: oData <= 16'h000a;
            14'h23fe: oData <= 16'h0000;
            14'h23ff: oData <= 16'h0000;
            14'h2400: oData <= 16'h0000;
            14'h2401: oData <= 16'h0000;
            14'h2402: oData <= 16'h0000;
            14'h2403: oData <= 16'h0000;
            14'h2404: oData <= 16'h0000;
            14'h2405: oData <= 16'h0000;
            14'h2406: oData <= 16'h0000;
            14'h2407: oData <= 16'ha800;
            14'h2408: oData <= 16'h0aaa;
            14'h2409: oData <= 16'h0000;
            14'h240a: oData <= 16'h0000;
            14'h240b: oData <= 16'haa00;
            14'h240c: oData <= 16'haaaa;
            14'h240d: oData <= 16'h0aaa;
            14'h240e: oData <= 16'haa80;
            14'h240f: oData <= 16'haaaa;
            14'h2410: oData <= 16'h2aaa;
            14'h2411: oData <= 16'h0000;
            14'h2412: oData <= 16'h0000;
            14'h2413: oData <= 16'h0000;
            14'h2414: oData <= 16'h0000;
            14'h2415: oData <= 16'h0000;
            14'h2416: oData <= 16'h0000;
            14'h2417: oData <= 16'h0000;
            14'h2418: oData <= 16'h0000;
            14'h2419: oData <= 16'h0000;
            14'h241a: oData <= 16'h0000;
            14'h241b: oData <= 16'h8000;
            14'h241c: oData <= 16'haaaa;
            14'h241d: oData <= 16'h0000;
            14'h241e: oData <= 16'h0000;
            14'h241f: oData <= 16'haa80;
            14'h2420: oData <= 16'haaaa;
            14'h2421: oData <= 16'haaaa;
            14'h2422: oData <= 16'haaaa;
            14'h2423: oData <= 16'haaaa;
            14'h2424: oData <= 16'h00aa;
            14'h2425: oData <= 16'h0000;
            14'h2426: oData <= 16'h0000;
            14'h2427: oData <= 16'h0000;
            14'h2428: oData <= 16'h0000;
            14'h2429: oData <= 16'h0000;
            14'h242a: oData <= 16'h0000;
            14'h242b: oData <= 16'h0000;
            14'h242c: oData <= 16'h0000;
            14'h242d: oData <= 16'h0000;
            14'h242e: oData <= 16'h0000;
            14'h242f: oData <= 16'h0000;
            14'h2430: oData <= 16'haaaa;
            14'h2431: oData <= 16'h0002;
            14'h2432: oData <= 16'h0000;
            14'h2433: oData <= 16'haaa0;
            14'h2434: oData <= 16'haaaa;
            14'h2435: oData <= 16'haaaa;
            14'h2436: oData <= 16'haaaa;
            14'h2437: oData <= 16'haaaa;
            14'h2438: oData <= 16'h0002;
            14'h2439: oData <= 16'h0000;
            14'h243a: oData <= 16'h0000;
            14'h243b: oData <= 16'h0000;
            14'h243c: oData <= 16'h0000;
            14'h243d: oData <= 16'h0000;
            14'h243e: oData <= 16'h0000;
            14'h243f: oData <= 16'h0000;
            14'h2440: oData <= 16'h0000;
            14'h2441: oData <= 16'h0000;
            14'h2442: oData <= 16'h0000;
            14'h2443: oData <= 16'h0000;
            14'h2444: oData <= 16'haaa0;
            14'h2445: oData <= 16'h0002;
            14'h2446: oData <= 16'h0000;
            14'h2447: oData <= 16'haaa8;
            14'h2448: oData <= 16'haaaa;
            14'h2449: oData <= 16'haaaa;
            14'h244a: oData <= 16'haaaa;
            14'h244b: oData <= 16'h0aaa;
            14'h244c: oData <= 16'h0000;
            14'h244d: oData <= 16'h0000;
            14'h244e: oData <= 16'h0000;
            14'h244f: oData <= 16'h0000;
            14'h2450: oData <= 16'h0000;
            14'h2451: oData <= 16'h0000;
            14'h2452: oData <= 16'h0000;
            14'h2453: oData <= 16'h0000;
            14'h2454: oData <= 16'h0000;
            14'h2455: oData <= 16'h0000;
            14'h2456: oData <= 16'h0000;
            14'h2457: oData <= 16'h0000;
            14'h2458: oData <= 16'haa00;
            14'h2459: oData <= 16'h0000;
            14'h245a: oData <= 16'h0000;
            14'h245b: oData <= 16'h0aaa;
            14'h245c: oData <= 16'ha000;
            14'h245d: oData <= 16'haaaa;
            14'h245e: oData <= 16'haaaa;
            14'h245f: oData <= 16'h002a;
            14'h2460: oData <= 16'h0000;
            14'h2461: oData <= 16'h0000;
            14'h2462: oData <= 16'h0000;
            14'h2463: oData <= 16'h0000;
            14'h2464: oData <= 16'h0000;
            14'h2465: oData <= 16'h0000;
            14'h2466: oData <= 16'h0000;
            14'h2467: oData <= 16'h0000;
            14'h2468: oData <= 16'h0000;
            14'h2469: oData <= 16'h0000;
            14'h246a: oData <= 16'h0000;
            14'h246b: oData <= 16'h0000;
            14'h246c: oData <= 16'h0000;
            14'h246d: oData <= 16'h0000;
            14'h246e: oData <= 16'h8000;
            14'h246f: oData <= 16'h02aa;
            14'h2470: oData <= 16'h0000;
            14'h2471: oData <= 16'ha800;
            14'h2472: oData <= 16'h2aaa;
            14'h2473: oData <= 16'h0000;
            14'h2474: oData <= 16'h0000;
            14'h2475: oData <= 16'h0000;
            14'h2476: oData <= 16'h0000;
            14'h2477: oData <= 16'h0000;
            14'h2478: oData <= 16'h0000;
            14'h2479: oData <= 16'h0000;
            14'h247a: oData <= 16'h0000;
            14'h247b: oData <= 16'h0000;
            14'h247c: oData <= 16'h0000;
            14'h247d: oData <= 16'h0000;
            14'h247e: oData <= 16'h0000;
            14'h247f: oData <= 16'h0000;
            14'h2480: oData <= 16'h0000;
            14'h2481: oData <= 16'h0000;
            14'h2482: oData <= 16'ha000;
            14'h2483: oData <= 16'h00aa;
            14'h2484: oData <= 16'h0000;
            14'h2485: oData <= 16'h0000;
            14'h2486: oData <= 16'h0000;
            14'h2487: oData <= 16'h0000;
            14'h2488: oData <= 16'h0000;
            14'h2489: oData <= 16'h0000;
            14'h248a: oData <= 16'h0000;
            14'h248b: oData <= 16'h0000;
            14'h248c: oData <= 16'h0000;
            14'h248d: oData <= 16'h0000;
            14'h248e: oData <= 16'h0000;
            14'h248f: oData <= 16'h0000;
            14'h2490: oData <= 16'h0000;
            14'h2491: oData <= 16'h0000;
            14'h2492: oData <= 16'h0000;
            14'h2493: oData <= 16'h0000;
            14'h2494: oData <= 16'h0000;
            14'h2495: oData <= 16'h0000;
            14'h2496: oData <= 16'ha800;
            14'h2497: oData <= 16'h002a;
            14'h2498: oData <= 16'h0000;
            14'h2499: oData <= 16'h0000;
            14'h249a: oData <= 16'h0000;
            14'h249b: oData <= 16'h0000;
            14'h249c: oData <= 16'h0000;
            14'h249d: oData <= 16'h0000;
            14'h249e: oData <= 16'h0000;
            14'h249f: oData <= 16'h0000;
            14'h24a0: oData <= 16'h0000;
            14'h24a1: oData <= 16'h0000;
            14'h24a2: oData <= 16'h0000;
            14'h24a3: oData <= 16'h0000;
            14'h24a4: oData <= 16'h0000;
            14'h24a5: oData <= 16'h0000;
            14'h24a6: oData <= 16'h0000;
            14'h24a7: oData <= 16'h0000;
            14'h24a8: oData <= 16'h0000;
            14'h24a9: oData <= 16'h0000;
            14'h24aa: oData <= 16'haa00;
            14'h24ab: oData <= 16'h000a;
            14'h24ac: oData <= 16'h0000;
            14'h24ad: oData <= 16'h0000;
            14'h24ae: oData <= 16'h0000;
            14'h24af: oData <= 16'h0000;
            14'h24b0: oData <= 16'h0000;
            14'h24b1: oData <= 16'h0000;
            14'h24b2: oData <= 16'h0000;
            14'h24b3: oData <= 16'h0000;
            14'h24b4: oData <= 16'h0000;
            14'h24b5: oData <= 16'h0000;
            14'h24b6: oData <= 16'h0000;
            14'h24b7: oData <= 16'h0000;
            14'h24b8: oData <= 16'h0000;
            14'h24b9: oData <= 16'h0000;
            14'h24ba: oData <= 16'h0000;
            14'h24bb: oData <= 16'h0000;
            14'h24bc: oData <= 16'h0000;
            14'h24bd: oData <= 16'h0000;
            14'h24be: oData <= 16'haa80;
            14'h24bf: oData <= 16'h0002;
            14'h24c0: oData <= 16'h0000;
            14'h24c1: oData <= 16'h0000;
            14'h24c2: oData <= 16'h0000;
            14'h24c3: oData <= 16'h0000;
            14'h24c4: oData <= 16'h0000;
            14'h24c5: oData <= 16'h0000;
            14'h24c6: oData <= 16'h0000;
            14'h24c7: oData <= 16'h0000;
            14'h24c8: oData <= 16'h0000;
            14'h24c9: oData <= 16'h0000;
            14'h24ca: oData <= 16'h0000;
            14'h24cb: oData <= 16'h0000;
            14'h24cc: oData <= 16'h0000;
            14'h24cd: oData <= 16'h0000;
            14'h24ce: oData <= 16'h0000;
            14'h24cf: oData <= 16'h0000;
            14'h24d0: oData <= 16'h0000;
            14'h24d1: oData <= 16'h0000;
            14'h24d2: oData <= 16'haaa8;
            14'h24d3: oData <= 16'h0000;
            14'h24d4: oData <= 16'h0000;
            14'h24d5: oData <= 16'h0000;
            14'h24d6: oData <= 16'h0000;
            14'h24d7: oData <= 16'h0000;
            14'h24d8: oData <= 16'h0000;
            14'h24d9: oData <= 16'h0000;
            14'h24da: oData <= 16'h0000;
            14'h24db: oData <= 16'h0000;
            14'h24dc: oData <= 16'h0000;
            14'h24dd: oData <= 16'h0000;
            14'h24de: oData <= 16'h0000;
            14'h24df: oData <= 16'h0000;
            14'h24e0: oData <= 16'h0000;
            14'h24e1: oData <= 16'h0000;
            14'h24e2: oData <= 16'h0000;
            14'h24e3: oData <= 16'h0000;
            14'h24e4: oData <= 16'h0000;
            14'h24e5: oData <= 16'h0000;
            14'h24e6: oData <= 16'h2aaa;
            14'h24e7: oData <= 16'h0000;
            14'h24e8: oData <= 16'h0000;
            14'h24e9: oData <= 16'h0000;
            14'h24ea: oData <= 16'h0000;
            14'h24eb: oData <= 16'h0000;
            14'h24ec: oData <= 16'h0000;
            14'h24ed: oData <= 16'h0000;
            14'h24ee: oData <= 16'h0000;
            14'h24ef: oData <= 16'h0000;
            14'h24f0: oData <= 16'h0000;
            14'h24f1: oData <= 16'h0000;
            14'h24f2: oData <= 16'h0000;
            14'h24f3: oData <= 16'h0000;
            14'h24f4: oData <= 16'h0000;
            14'h24f5: oData <= 16'h0000;
            14'h24f6: oData <= 16'h0000;
            14'h24f7: oData <= 16'h0000;
            14'h24f8: oData <= 16'h0000;
            14'h24f9: oData <= 16'h0000;
            14'h24fa: oData <= 16'h0aaa;
            14'h24fb: oData <= 16'h0000;
            14'h24fc: oData <= 16'h0000;
            14'h24fd: oData <= 16'h0000;
            14'h24fe: oData <= 16'h0000;
            14'h24ff: oData <= 16'h0000;
            14'h2500: oData <= 16'h0000;
            14'h2501: oData <= 16'h0000;
            14'h2502: oData <= 16'h0000;
            14'h2503: oData <= 16'h0000;
            14'h2504: oData <= 16'h0000;
            14'h2505: oData <= 16'h0000;
            14'h2506: oData <= 16'h0000;
            14'h2507: oData <= 16'h0000;
            14'h2508: oData <= 16'h0000;
            14'h2509: oData <= 16'h0000;
            14'h250a: oData <= 16'h0000;
            14'h250b: oData <= 16'h0000;
            14'h250c: oData <= 16'h0000;
            14'h250d: oData <= 16'h0000;
            14'h250e: oData <= 16'h02aa;
            14'h250f: oData <= 16'h0000;
            14'h2510: oData <= 16'h0000;
            14'h2511: oData <= 16'h0000;
            14'h2512: oData <= 16'h0000;
            14'h2513: oData <= 16'h0000;
            14'h2514: oData <= 16'h0000;
            14'h2515: oData <= 16'h0000;
            14'h2516: oData <= 16'h0000;
            14'h2517: oData <= 16'h0000;
            14'h2518: oData <= 16'h0000;
            14'h2519: oData <= 16'h0000;
            14'h251a: oData <= 16'h0000;
            14'h251b: oData <= 16'h0000;
            14'h251c: oData <= 16'h0000;
            14'h251d: oData <= 16'h0000;
            14'h251e: oData <= 16'h0000;
            14'h251f: oData <= 16'h0000;
            14'h2520: oData <= 16'h0000;
            14'h2521: oData <= 16'h0000;
            14'h2522: oData <= 16'h00a8;
            14'h2523: oData <= 16'h0000;
            14'h2524: oData <= 16'h0000;
            14'h2525: oData <= 16'h0000;
            14'h2526: oData <= 16'h0000;
            14'h2527: oData <= 16'h0000;
            14'h2528: oData <= 16'h0000;
            14'h2529: oData <= 16'h0000;
            14'h252a: oData <= 16'h0000;
            14'h252b: oData <= 16'h0000;
            14'h252c: oData <= 16'h0000;
            14'h252d: oData <= 16'h0000;
            14'h252e: oData <= 16'h0000;
            14'h252f: oData <= 16'h0000;
            14'h2530: oData <= 16'h0000;
            14'h2531: oData <= 16'h0000;
            14'h2532: oData <= 16'h0000;
            14'h2533: oData <= 16'h0000;
            14'h2534: oData <= 16'h0000;
            14'h2535: oData <= 16'h0000;
            14'h2536: oData <= 16'h0000;
            14'h2537: oData <= 16'h0000;
            14'h2538: oData <= 16'h0000;
            14'h2539: oData <= 16'h0000;
            14'h253a: oData <= 16'h0000;
            14'h253b: oData <= 16'h0000;
            14'h253c: oData <= 16'h0000;
            14'h253d: oData <= 16'h0000;
            14'h253e: oData <= 16'h0000;
            14'h253f: oData <= 16'h0000;
            14'h2540: oData <= 16'h0000;
            14'h2541: oData <= 16'h0000;
            14'h2542: oData <= 16'h0000;
            14'h2543: oData <= 16'h0000;
            14'h2544: oData <= 16'h0000;
            14'h2545: oData <= 16'h0000;
            14'h2546: oData <= 16'h0000;
            14'h2547: oData <= 16'h0000;
            14'h2548: oData <= 16'h0000;
            14'h2549: oData <= 16'h0000;
            14'h254a: oData <= 16'h0000;
            14'h254b: oData <= 16'h0000;
            14'h254c: oData <= 16'h0000;
            14'h254d: oData <= 16'h0000;
            14'h254e: oData <= 16'h0000;
            14'h254f: oData <= 16'h0000;
            14'h2550: oData <= 16'h0000;
            14'h2551: oData <= 16'h0000;
            14'h2552: oData <= 16'h0000;
            14'h2553: oData <= 16'h0000;
            14'h2554: oData <= 16'h0000;
            14'h2555: oData <= 16'h0000;
            14'h2556: oData <= 16'h0000;
            14'h2557: oData <= 16'h0000;
            14'h2558: oData <= 16'h0000;
            14'h2559: oData <= 16'h0000;
            14'h255a: oData <= 16'h0000;
            14'h255b: oData <= 16'h0000;
            14'h255c: oData <= 16'h0000;
            14'h255d: oData <= 16'h0000;
            14'h255e: oData <= 16'h0000;
            14'h255f: oData <= 16'h0000;
            14'h2560: oData <= 16'h0000;
            14'h2561: oData <= 16'h0000;
            14'h2562: oData <= 16'h0000;
            14'h2563: oData <= 16'h0000;
            14'h2564: oData <= 16'h0000;
            14'h2565: oData <= 16'h0000;
            14'h2566: oData <= 16'h0000;
            14'h2567: oData <= 16'h0000;
            14'h2568: oData <= 16'h0000;
            14'h2569: oData <= 16'h0000;
            14'h256a: oData <= 16'h0000;
            14'h256b: oData <= 16'h0000;
            14'h256c: oData <= 16'h0000;
            14'h256d: oData <= 16'h0000;
            14'h256e: oData <= 16'h0000;
            14'h256f: oData <= 16'h0000;
            14'h2570: oData <= 16'h0000;
            14'h2571: oData <= 16'h0000;
            14'h2572: oData <= 16'h0000;
            14'h2573: oData <= 16'h0000;
            14'h2574: oData <= 16'h0000;
            14'h2575: oData <= 16'h0000;
            14'h2576: oData <= 16'h0000;
            14'h2577: oData <= 16'h0000;
            14'h2578: oData <= 16'h0000;
            14'h2579: oData <= 16'h0000;
            14'h257a: oData <= 16'h0000;
            14'h257b: oData <= 16'h0000;
            14'h257c: oData <= 16'h0000;
            14'h257d: oData <= 16'h0000;
            14'h257e: oData <= 16'h0000;
            14'h257f: oData <= 16'h0000;
            14'h2580: oData <= 16'h0000;
            14'h2581: oData <= 16'h0000;
            14'h2582: oData <= 16'h0000;
            14'h2583: oData <= 16'h0000;
            14'h2584: oData <= 16'h0000;
            14'h2585: oData <= 16'h0000;
            14'h2586: oData <= 16'h0000;
            14'h2587: oData <= 16'h0000;
            14'h2588: oData <= 16'h0000;
            14'h2589: oData <= 16'h0000;
            14'h258a: oData <= 16'h0000;
            14'h258b: oData <= 16'h0000;
            14'h258c: oData <= 16'h0000;
            14'h258d: oData <= 16'h0000;
            14'h258e: oData <= 16'h0000;
            14'h258f: oData <= 16'h0000;
            14'h2590: oData <= 16'h0000;
            14'h2591: oData <= 16'h0000;
            14'h2592: oData <= 16'h0000;
            14'h2593: oData <= 16'h0000;
            14'h2594: oData <= 16'h0000;
            14'h2595: oData <= 16'h0000;
            14'h2596: oData <= 16'h0000;
            14'h2597: oData <= 16'h0000;
            14'h2598: oData <= 16'h0000;
            14'h2599: oData <= 16'h0000;
            14'h259a: oData <= 16'h0000;
            14'h259b: oData <= 16'h0000;
            14'h259c: oData <= 16'h0000;
            14'h259d: oData <= 16'h0000;
            14'h259e: oData <= 16'h0000;
            14'h259f: oData <= 16'h0000;
            14'h25a0: oData <= 16'h0000;
            14'h25a1: oData <= 16'h0000;
            14'h25a2: oData <= 16'h0000;
            14'h25a3: oData <= 16'h0000;
            14'h25a4: oData <= 16'h0000;
            14'h25a5: oData <= 16'h0000;
            14'h25a6: oData <= 16'h0000;
            14'h25a7: oData <= 16'h0000;
            14'h25a8: oData <= 16'h0000;
            14'h25a9: oData <= 16'h0000;
            14'h25aa: oData <= 16'h0000;
            14'h25ab: oData <= 16'h0000;
            14'h25ac: oData <= 16'h0000;
            14'h25ad: oData <= 16'h0000;
            14'h25ae: oData <= 16'h0000;
            14'h25af: oData <= 16'h0000;
            14'h25b0: oData <= 16'h0000;
            14'h25b1: oData <= 16'h0000;
            14'h25b2: oData <= 16'h0000;
            14'h25b3: oData <= 16'h0000;
            14'h25b4: oData <= 16'h0000;
            14'h25b5: oData <= 16'h0000;
            14'h25b6: oData <= 16'h0000;
            14'h25b7: oData <= 16'h0000;
            14'h25b8: oData <= 16'h0000;
            14'h25b9: oData <= 16'h0000;
            14'h25ba: oData <= 16'h0000;
            14'h25bb: oData <= 16'h0000;
            14'h25bc: oData <= 16'h0000;
            14'h25bd: oData <= 16'h0000;
            14'h25be: oData <= 16'h0000;
            14'h25bf: oData <= 16'h0000;
            14'h25c0: oData <= 16'h0000;
            14'h25c1: oData <= 16'h0000;
            14'h25c2: oData <= 16'h0000;
            14'h25c3: oData <= 16'h0000;
            14'h25c4: oData <= 16'h0000;
            14'h25c5: oData <= 16'h0000;
            14'h25c6: oData <= 16'h0000;
            14'h25c7: oData <= 16'h0000;
            14'h25c8: oData <= 16'h0000;
            14'h25c9: oData <= 16'h0000;
            14'h25ca: oData <= 16'h0000;
            14'h25cb: oData <= 16'h0000;
            14'h25cc: oData <= 16'h0000;
            14'h25cd: oData <= 16'h0000;
            14'h25ce: oData <= 16'h0000;
            14'h25cf: oData <= 16'h0000;
            14'h25d0: oData <= 16'h0000;
            14'h25d1: oData <= 16'h0000;
            14'h25d2: oData <= 16'h0000;
            14'h25d3: oData <= 16'h0000;
            14'h25d4: oData <= 16'h0000;
            14'h25d5: oData <= 16'h0000;
            14'h25d6: oData <= 16'h0000;
            14'h25d7: oData <= 16'h0000;
            14'h25d8: oData <= 16'h0000;
            14'h25d9: oData <= 16'h0000;
            14'h25da: oData <= 16'h0000;
            14'h25db: oData <= 16'h0000;
            14'h25dc: oData <= 16'h0000;
            14'h25dd: oData <= 16'h0000;
            14'h25de: oData <= 16'h0000;
            14'h25df: oData <= 16'h0000;
            14'h25e0: oData <= 16'h0000;
            14'h25e1: oData <= 16'h0000;
            14'h25e2: oData <= 16'h0000;
            14'h25e3: oData <= 16'h0000;
            14'h25e4: oData <= 16'h0000;
            14'h25e5: oData <= 16'h0000;
            14'h25e6: oData <= 16'h0000;
            14'h25e7: oData <= 16'h0000;
            14'h25e8: oData <= 16'h0000;
            14'h25e9: oData <= 16'h0000;
            14'h25ea: oData <= 16'h0000;
            14'h25eb: oData <= 16'h0000;
            14'h25ec: oData <= 16'h0000;
            14'h25ed: oData <= 16'h0000;
            14'h25ee: oData <= 16'h0000;
            14'h25ef: oData <= 16'h0000;
            14'h25f0: oData <= 16'h0000;
            14'h25f1: oData <= 16'h0000;
            14'h25f2: oData <= 16'h0000;
            14'h25f3: oData <= 16'h0000;
            14'h25f4: oData <= 16'h0000;
            14'h25f5: oData <= 16'h0000;
            14'h25f6: oData <= 16'h0000;
            14'h25f7: oData <= 16'h0000;
            14'h25f8: oData <= 16'h0000;
            14'h25f9: oData <= 16'h0000;
            14'h25fa: oData <= 16'h0000;
            14'h25fb: oData <= 16'h0000;
            14'h25fc: oData <= 16'h0000;
            14'h25fd: oData <= 16'h0000;
            14'h25fe: oData <= 16'h0000;
            14'h25ff: oData <= 16'h0000;
            14'h2600: oData <= 16'h0000;
            14'h2601: oData <= 16'h0000;
            14'h2602: oData <= 16'h0000;
            14'h2603: oData <= 16'h0000;
            14'h2604: oData <= 16'h0000;
            14'h2605: oData <= 16'h0000;
            14'h2606: oData <= 16'h0000;
            14'h2607: oData <= 16'h0000;
            14'h2608: oData <= 16'h0000;
            14'h2609: oData <= 16'h0000;
            14'h260a: oData <= 16'h0000;
            14'h260b: oData <= 16'h0000;
            14'h260c: oData <= 16'h0000;
            14'h260d: oData <= 16'h0000;
            14'h260e: oData <= 16'h0000;
            14'h260f: oData <= 16'h0000;
            14'h2610: oData <= 16'h0000;
            14'h2611: oData <= 16'h0000;
            14'h2612: oData <= 16'h0000;
            14'h2613: oData <= 16'h0000;
            14'h2614: oData <= 16'h0000;
            14'h2615: oData <= 16'h0000;
            14'h2616: oData <= 16'h0000;
            14'h2617: oData <= 16'h0000;
            14'h2618: oData <= 16'h0000;
            14'h2619: oData <= 16'h0000;
            14'h261a: oData <= 16'h0000;
            14'h261b: oData <= 16'h0000;
            14'h261c: oData <= 16'h0000;
            14'h261d: oData <= 16'h0000;
            14'h261e: oData <= 16'h0000;
            14'h261f: oData <= 16'h0000;
            14'h2620: oData <= 16'h0000;
            14'h2621: oData <= 16'h0000;
            14'h2622: oData <= 16'h0000;
            14'h2623: oData <= 16'h0000;
            14'h2624: oData <= 16'h0000;
            14'h2625: oData <= 16'h0000;
            14'h2626: oData <= 16'h0000;
            14'h2627: oData <= 16'h0000;
            14'h2628: oData <= 16'h0000;
            14'h2629: oData <= 16'h0000;
            14'h262a: oData <= 16'h0000;
            14'h262b: oData <= 16'h0000;
            14'h262c: oData <= 16'h0000;
            14'h262d: oData <= 16'h0000;
            14'h262e: oData <= 16'h0000;
            14'h262f: oData <= 16'h0000;
            14'h2630: oData <= 16'h0000;
            14'h2631: oData <= 16'h0000;
            14'h2632: oData <= 16'h0000;
            14'h2633: oData <= 16'h0000;
            14'h2634: oData <= 16'h0000;
            14'h2635: oData <= 16'h0000;
            14'h2636: oData <= 16'h0000;
            14'h2637: oData <= 16'h0000;
            14'h2638: oData <= 16'h0000;
            14'h2639: oData <= 16'h0000;
            14'h263a: oData <= 16'h0000;
            14'h263b: oData <= 16'h0000;
            14'h263c: oData <= 16'h0000;
            14'h263d: oData <= 16'h0000;
            14'h263e: oData <= 16'h0000;
            14'h263f: oData <= 16'h0000;
            14'h2640: oData <= 16'h0000;
            14'h2641: oData <= 16'h0000;
            14'h2642: oData <= 16'h0000;
            14'h2643: oData <= 16'h0000;
            14'h2644: oData <= 16'h0000;
            14'h2645: oData <= 16'h0000;
            14'h2646: oData <= 16'h0000;
            14'h2647: oData <= 16'h0000;
            14'h2648: oData <= 16'h0000;
            14'h2649: oData <= 16'h0000;
            14'h264a: oData <= 16'h0000;
            14'h264b: oData <= 16'h0000;
            14'h264c: oData <= 16'h0000;
            14'h264d: oData <= 16'h0000;
            14'h264e: oData <= 16'h0000;
            14'h264f: oData <= 16'h0000;
            14'h2650: oData <= 16'h0000;
            14'h2651: oData <= 16'h0000;
            14'h2652: oData <= 16'h0000;
            14'h2653: oData <= 16'h0000;
            14'h2654: oData <= 16'h0000;
            14'h2655: oData <= 16'h0000;
            14'h2656: oData <= 16'h0000;
            14'h2657: oData <= 16'h0000;
            14'h2658: oData <= 16'h0000;
            14'h2659: oData <= 16'h0000;
            14'h265a: oData <= 16'h0000;
            14'h265b: oData <= 16'h0000;
            14'h265c: oData <= 16'h0000;
            14'h265d: oData <= 16'h0000;
            14'h265e: oData <= 16'h0000;
            14'h265f: oData <= 16'h0000;
            14'h2660: oData <= 16'h0000;
            14'h2661: oData <= 16'h0000;
            14'h2662: oData <= 16'h0000;
            14'h2663: oData <= 16'h0000;
            14'h2664: oData <= 16'h0000;
            14'h2665: oData <= 16'h0000;
            14'h2666: oData <= 16'h0000;
            14'h2667: oData <= 16'h0000;
            14'h2668: oData <= 16'h0000;
            14'h2669: oData <= 16'h0000;
            14'h266a: oData <= 16'h0000;
            14'h266b: oData <= 16'h0000;
            14'h266c: oData <= 16'h0000;
            14'h266d: oData <= 16'h0000;
            14'h266e: oData <= 16'h0000;
            14'h266f: oData <= 16'h0000;
            14'h2670: oData <= 16'h0000;
            14'h2671: oData <= 16'h0000;
            14'h2672: oData <= 16'h0000;
            14'h2673: oData <= 16'h0000;
            14'h2674: oData <= 16'h0000;
            14'h2675: oData <= 16'h0000;
            14'h2676: oData <= 16'h0000;
            14'h2677: oData <= 16'h0000;
            14'h2678: oData <= 16'h0000;
            14'h2679: oData <= 16'h0000;
            14'h267a: oData <= 16'h0000;
            14'h267b: oData <= 16'h0000;
            14'h267c: oData <= 16'h0000;
            14'h267d: oData <= 16'h0000;
            14'h267e: oData <= 16'h0000;
            14'h267f: oData <= 16'h0000;
            14'h2680: oData <= 16'h0000;
            14'h2681: oData <= 16'h0000;
            14'h2682: oData <= 16'h0000;
            14'h2683: oData <= 16'h0000;
            14'h2684: oData <= 16'h0000;
            14'h2685: oData <= 16'h0000;
            14'h2686: oData <= 16'h0000;
            14'h2687: oData <= 16'h0000;
            14'h2688: oData <= 16'h0000;
            14'h2689: oData <= 16'h0000;
            14'h268a: oData <= 16'h0000;
            14'h268b: oData <= 16'h0000;
            14'h268c: oData <= 16'h0000;
            14'h268d: oData <= 16'h0000;
            14'h268e: oData <= 16'h0000;
            14'h268f: oData <= 16'h0000;
            14'h2690: oData <= 16'h0000;
            14'h2691: oData <= 16'h0000;
            14'h2692: oData <= 16'h0000;
            14'h2693: oData <= 16'h0000;
            14'h2694: oData <= 16'h0000;
            14'h2695: oData <= 16'h0000;
            14'h2696: oData <= 16'h0000;
            14'h2697: oData <= 16'h0000;
            14'h2698: oData <= 16'h0000;
            14'h2699: oData <= 16'h0000;
            14'h269a: oData <= 16'h0000;
            14'h269b: oData <= 16'h0000;
            14'h269c: oData <= 16'h0000;
            14'h269d: oData <= 16'h0000;
            14'h269e: oData <= 16'h0000;
            14'h269f: oData <= 16'h0000;
            14'h26a0: oData <= 16'h0000;
            14'h26a1: oData <= 16'h0000;
            14'h26a2: oData <= 16'h0000;
            14'h26a3: oData <= 16'h0000;
            14'h26a4: oData <= 16'h0000;
            14'h26a5: oData <= 16'h0000;
            14'h26a6: oData <= 16'h0000;
            14'h26a7: oData <= 16'h0000;
            14'h26a8: oData <= 16'h0000;
            14'h26a9: oData <= 16'h0000;
            14'h26aa: oData <= 16'h0000;
            14'h26ab: oData <= 16'h0000;
            14'h26ac: oData <= 16'h0000;
            14'h26ad: oData <= 16'h0000;
            14'h26ae: oData <= 16'h0000;
            14'h26af: oData <= 16'h0000;
            14'h26b0: oData <= 16'h0000;
            14'h26b1: oData <= 16'h0000;
            14'h26b2: oData <= 16'h0000;
            14'h26b3: oData <= 16'h0000;
            14'h26b4: oData <= 16'h0000;
            14'h26b5: oData <= 16'h0000;
            14'h26b6: oData <= 16'h0000;
            14'h26b7: oData <= 16'h0000;
            14'h26b8: oData <= 16'h0000;
            14'h26b9: oData <= 16'h0000;
            14'h26ba: oData <= 16'h0000;
            14'h26bb: oData <= 16'h0000;
            14'h26bc: oData <= 16'h0000;
            14'h26bd: oData <= 16'h0000;
            14'h26be: oData <= 16'h0000;
            14'h26bf: oData <= 16'h0000;
            14'h26c0: oData <= 16'h0000;
            14'h26c1: oData <= 16'h0000;
            14'h26c2: oData <= 16'h0000;
            14'h26c3: oData <= 16'h0000;
            14'h26c4: oData <= 16'h0000;
            14'h26c5: oData <= 16'h0000;
            14'h26c6: oData <= 16'h0000;
            14'h26c7: oData <= 16'h0000;
            14'h26c8: oData <= 16'h0000;
            14'h26c9: oData <= 16'h0000;
            14'h26ca: oData <= 16'h0000;
            14'h26cb: oData <= 16'h0000;
            14'h26cc: oData <= 16'h0000;
            14'h26cd: oData <= 16'h0000;
            14'h26ce: oData <= 16'h0000;
            14'h26cf: oData <= 16'h0000;
            14'h26d0: oData <= 16'h0000;
            14'h26d1: oData <= 16'h0000;
            14'h26d2: oData <= 16'h0000;
            14'h26d3: oData <= 16'h0000;
            14'h26d4: oData <= 16'h0000;
            14'h26d5: oData <= 16'h0000;
            14'h26d6: oData <= 16'h0000;
            14'h26d7: oData <= 16'h0000;
            14'h26d8: oData <= 16'h0000;
            14'h26d9: oData <= 16'h0000;
            14'h26da: oData <= 16'h0000;
            14'h26db: oData <= 16'h0000;
            14'h26dc: oData <= 16'h0000;
            14'h26dd: oData <= 16'h0000;
            14'h26de: oData <= 16'h0000;
            14'h26df: oData <= 16'h0000;
            14'h26e0: oData <= 16'h0000;
            14'h26e1: oData <= 16'h0000;
            14'h26e2: oData <= 16'h0000;
            14'h26e3: oData <= 16'h0000;
            14'h26e4: oData <= 16'h0000;
            14'h26e5: oData <= 16'h0000;
            14'h26e6: oData <= 16'h0000;
            14'h26e7: oData <= 16'h0000;
            14'h26e8: oData <= 16'h0000;
            14'h26e9: oData <= 16'h0000;
            14'h26ea: oData <= 16'h0000;
            14'h26eb: oData <= 16'h0000;
            14'h26ec: oData <= 16'h0000;
            14'h26ed: oData <= 16'h0000;
            14'h26ee: oData <= 16'h0000;
            14'h26ef: oData <= 16'h0000;
            14'h26f0: oData <= 16'h0000;
            14'h26f1: oData <= 16'h0000;
            14'h26f2: oData <= 16'h0000;
            14'h26f3: oData <= 16'h0000;
            14'h26f4: oData <= 16'h0000;
            14'h26f5: oData <= 16'h0000;
            14'h26f6: oData <= 16'h0000;
            14'h26f7: oData <= 16'h0000;
            14'h26f8: oData <= 16'h0000;
            14'h26f9: oData <= 16'h0000;
            14'h26fa: oData <= 16'h0000;
            14'h26fb: oData <= 16'h0000;
            14'h26fc: oData <= 16'h0000;
            14'h26fd: oData <= 16'h0000;
            14'h26fe: oData <= 16'h0000;
            14'h26ff: oData <= 16'h0000;
            14'h2700: oData <= 16'h0000;
            14'h2701: oData <= 16'h0000;
            14'h2702: oData <= 16'h0000;
            14'h2703: oData <= 16'h0000;
            14'h2704: oData <= 16'h0000;
            14'h2705: oData <= 16'h0000;
            14'h2706: oData <= 16'h0000;
            14'h2707: oData <= 16'h0000;
            14'h2708: oData <= 16'h0000;
            14'h2709: oData <= 16'h0000;
            14'h270a: oData <= 16'h0000;
            14'h270b: oData <= 16'h0000;
            14'h270c: oData <= 16'h0000;
            14'h270d: oData <= 16'h0000;
            14'h270e: oData <= 16'h0000;
            14'h270f: oData <= 16'h0000;
            14'h2710: oData <= 16'h0000;
            14'h2711: oData <= 16'h0000;
            14'h2712: oData <= 16'h0000;
            14'h2713: oData <= 16'h0000;
            14'h2714: oData <= 16'h0000;
            14'h2715: oData <= 16'h0000;
            14'h2716: oData <= 16'h0000;
            14'h2717: oData <= 16'h0000;
            14'h2718: oData <= 16'h0000;
            14'h2719: oData <= 16'h0000;
            14'h271a: oData <= 16'h0000;
            14'h271b: oData <= 16'h0000;
            14'h271c: oData <= 16'h0000;
            14'h271d: oData <= 16'h0000;
            14'h271e: oData <= 16'h0000;
            14'h271f: oData <= 16'h0000;
            14'h2720: oData <= 16'h0000;
            14'h2721: oData <= 16'h0000;
            14'h2722: oData <= 16'h0000;
            14'h2723: oData <= 16'h0000;
            14'h2724: oData <= 16'h0000;
            14'h2725: oData <= 16'h0000;
            14'h2726: oData <= 16'h0000;
            14'h2727: oData <= 16'h0000;
            14'h2728: oData <= 16'h0000;
            14'h2729: oData <= 16'h0000;
            14'h272a: oData <= 16'h0000;
            14'h272b: oData <= 16'h0000;
            14'h272c: oData <= 16'h0000;
            14'h272d: oData <= 16'h0000;
            14'h272e: oData <= 16'h0000;
            14'h272f: oData <= 16'h0000;
            14'h2730: oData <= 16'h0000;
            14'h2731: oData <= 16'h0000;
            14'h2732: oData <= 16'h0000;
            14'h2733: oData <= 16'h0000;
            14'h2734: oData <= 16'h0000;
            14'h2735: oData <= 16'h0000;
            14'h2736: oData <= 16'h0000;
            14'h2737: oData <= 16'h0000;
            14'h2738: oData <= 16'h0000;
            14'h2739: oData <= 16'h0000;
            14'h273a: oData <= 16'h0000;
            14'h273b: oData <= 16'h0000;
            14'h273c: oData <= 16'h0000;
            14'h273d: oData <= 16'h0000;
            14'h273e: oData <= 16'h0000;
            14'h273f: oData <= 16'h0000;
            14'h2740: oData <= 16'h0000;
            14'h2741: oData <= 16'h0000;
            14'h2742: oData <= 16'h0000;
            14'h2743: oData <= 16'h0000;
            14'h2744: oData <= 16'h0000;
            14'h2745: oData <= 16'h0000;
            14'h2746: oData <= 16'h0000;
            14'h2747: oData <= 16'h0000;
            14'h2748: oData <= 16'h0000;
            14'h2749: oData <= 16'h0000;
            14'h274a: oData <= 16'h0000;
            14'h274b: oData <= 16'h0000;
            14'h274c: oData <= 16'h0000;
            14'h274d: oData <= 16'h0000;
            14'h274e: oData <= 16'h0000;
            14'h274f: oData <= 16'h0000;
            14'h2750: oData <= 16'h0000;
            14'h2751: oData <= 16'h0000;
            14'h2752: oData <= 16'h0000;
            14'h2753: oData <= 16'h0000;
            14'h2754: oData <= 16'h0000;
            14'h2755: oData <= 16'h0000;
            14'h2756: oData <= 16'h0000;
            14'h2757: oData <= 16'h0000;
            14'h2758: oData <= 16'h0000;
            14'h2759: oData <= 16'h0000;
            14'h275a: oData <= 16'h0000;
            14'h275b: oData <= 16'h0000;
            14'h275c: oData <= 16'h0000;
            14'h275d: oData <= 16'h0000;
            14'h275e: oData <= 16'h0000;
            14'h275f: oData <= 16'h0000;
            14'h2760: oData <= 16'h0000;
            14'h2761: oData <= 16'h0000;
            14'h2762: oData <= 16'h0000;
            14'h2763: oData <= 16'h0000;
            14'h2764: oData <= 16'h0000;
            14'h2765: oData <= 16'h0000;
            14'h2766: oData <= 16'h0000;
            14'h2767: oData <= 16'h0000;
            14'h2768: oData <= 16'h0000;
            14'h2769: oData <= 16'h0000;
            14'h276a: oData <= 16'h0000;
            14'h276b: oData <= 16'h0000;
            14'h276c: oData <= 16'h0000;
            14'h276d: oData <= 16'h0000;
            14'h276e: oData <= 16'h0000;
            14'h276f: oData <= 16'h0000;
            14'h2770: oData <= 16'h0000;
            14'h2771: oData <= 16'h0000;
            14'h2772: oData <= 16'h0000;
            14'h2773: oData <= 16'h0000;
            14'h2774: oData <= 16'h0000;
            14'h2775: oData <= 16'h0000;
            14'h2776: oData <= 16'h0000;
            14'h2777: oData <= 16'h0000;
            14'h2778: oData <= 16'h0000;
            14'h2779: oData <= 16'h0000;
            14'h277a: oData <= 16'h0000;
            14'h277b: oData <= 16'h0000;
            14'h277c: oData <= 16'h0000;
            14'h277d: oData <= 16'h0000;
            14'h277e: oData <= 16'h0000;
            14'h277f: oData <= 16'h0000;
            14'h2780: oData <= 16'h0000;
            14'h2781: oData <= 16'h0000;
            14'h2782: oData <= 16'h0000;
            14'h2783: oData <= 16'h0000;
            14'h2784: oData <= 16'h0000;
            14'h2785: oData <= 16'h0000;
            14'h2786: oData <= 16'h0000;
            14'h2787: oData <= 16'h0000;
            14'h2788: oData <= 16'h0000;
            14'h2789: oData <= 16'h0000;
            14'h278a: oData <= 16'h0000;
            14'h278b: oData <= 16'h0000;
            14'h278c: oData <= 16'h0000;
            14'h278d: oData <= 16'h0000;
            14'h278e: oData <= 16'h0000;
            14'h278f: oData <= 16'h0000;
            14'h2790: oData <= 16'h0000;
            14'h2791: oData <= 16'h0000;
            14'h2792: oData <= 16'h0000;
            14'h2793: oData <= 16'h0000;
            14'h2794: oData <= 16'h0000;
            14'h2795: oData <= 16'h0000;
            14'h2796: oData <= 16'h0000;
            14'h2797: oData <= 16'h0000;
            14'h2798: oData <= 16'h0000;
            14'h2799: oData <= 16'h0000;
            14'h279a: oData <= 16'h0000;
            14'h279b: oData <= 16'h0000;
            14'h279c: oData <= 16'h0000;
            14'h279d: oData <= 16'h0000;
            14'h279e: oData <= 16'h0000;
            14'h279f: oData <= 16'h0000;
            14'h27a0: oData <= 16'h0000;
            14'h27a1: oData <= 16'h0000;
            14'h27a2: oData <= 16'h0000;
            14'h27a3: oData <= 16'h0000;
            14'h27a4: oData <= 16'h0000;
            14'h27a5: oData <= 16'h0000;
            14'h27a6: oData <= 16'h0000;
            14'h27a7: oData <= 16'h0000;
            14'h27a8: oData <= 16'h0000;
            14'h27a9: oData <= 16'h0000;
            14'h27aa: oData <= 16'h0000;
            14'h27ab: oData <= 16'h0000;
            14'h27ac: oData <= 16'h0000;
            14'h27ad: oData <= 16'h0000;
            14'h27ae: oData <= 16'h0000;
            14'h27af: oData <= 16'h0000;
            14'h27b0: oData <= 16'h0000;
            14'h27b1: oData <= 16'h0000;
            14'h27b2: oData <= 16'h0000;
            14'h27b3: oData <= 16'h0000;
            14'h27b4: oData <= 16'h0000;
            14'h27b5: oData <= 16'h0000;
            14'h27b6: oData <= 16'h0000;
            14'h27b7: oData <= 16'h0000;
            14'h27b8: oData <= 16'h0000;
            14'h27b9: oData <= 16'h0000;
            14'h27ba: oData <= 16'h0000;
            14'h27bb: oData <= 16'h0000;
            14'h27bc: oData <= 16'h0000;
            14'h27bd: oData <= 16'h0000;
            14'h27be: oData <= 16'h0000;
            14'h27bf: oData <= 16'h0000;
            14'h27c0: oData <= 16'h0000;
            14'h27c1: oData <= 16'h0000;
            14'h27c2: oData <= 16'h0000;
            14'h27c3: oData <= 16'h0000;
            14'h27c4: oData <= 16'h0000;
            14'h27c5: oData <= 16'h0000;
            14'h27c6: oData <= 16'h0000;
            14'h27c7: oData <= 16'h0000;
            14'h27c8: oData <= 16'h0000;
            14'h27c9: oData <= 16'h0000;
            14'h27ca: oData <= 16'h0000;
            14'h27cb: oData <= 16'h0000;
            14'h27cc: oData <= 16'h0000;
            14'h27cd: oData <= 16'h0000;
            14'h27ce: oData <= 16'h0000;
            14'h27cf: oData <= 16'h0000;
            14'h27d0: oData <= 16'h0000;
            14'h27d1: oData <= 16'h0000;
            14'h27d2: oData <= 16'h0000;
            14'h27d3: oData <= 16'h0000;
            14'h27d4: oData <= 16'h0000;
            14'h27d5: oData <= 16'h0000;
            14'h27d6: oData <= 16'h0000;
            14'h27d7: oData <= 16'h0000;
            14'h27d8: oData <= 16'h0000;
            14'h27d9: oData <= 16'h0000;
            14'h27da: oData <= 16'h0000;
            14'h27db: oData <= 16'h0000;
            14'h27dc: oData <= 16'h0000;
            14'h27dd: oData <= 16'h0000;
            14'h27de: oData <= 16'h0000;
            14'h27df: oData <= 16'h0000;
            14'h27e0: oData <= 16'h0000;
            14'h27e1: oData <= 16'h0000;
            14'h27e2: oData <= 16'h0000;
            14'h27e3: oData <= 16'h0000;
            14'h27e4: oData <= 16'h0000;
            14'h27e5: oData <= 16'h0000;
            14'h27e6: oData <= 16'h0000;
            14'h27e7: oData <= 16'h0000;
            14'h27e8: oData <= 16'h0000;
            14'h27e9: oData <= 16'h0000;
            14'h27ea: oData <= 16'h0000;
            14'h27eb: oData <= 16'h0000;
            14'h27ec: oData <= 16'h0000;
            14'h27ed: oData <= 16'h0000;
            14'h27ee: oData <= 16'h0000;
            14'h27ef: oData <= 16'h0000;
            14'h27f0: oData <= 16'h0000;
            14'h27f1: oData <= 16'h0000;
            14'h27f2: oData <= 16'h0000;
            14'h27f3: oData <= 16'h0000;
            14'h27f4: oData <= 16'h0000;
            14'h27f5: oData <= 16'h0000;
            14'h27f6: oData <= 16'h0000;
            14'h27f7: oData <= 16'h0000;
            14'h27f8: oData <= 16'h0000;
            14'h27f9: oData <= 16'h0000;
            14'h27fa: oData <= 16'h0000;
            14'h27fb: oData <= 16'h0000;
            14'h27fc: oData <= 16'h0000;
            14'h27fd: oData <= 16'h0000;
            14'h27fe: oData <= 16'h0000;
            14'h27ff: oData <= 16'h0000;
            14'h2800: oData <= 16'h0000;
            14'h2801: oData <= 16'h0000;
            14'h2802: oData <= 16'h0000;
            14'h2803: oData <= 16'h0000;
            14'h2804: oData <= 16'h0000;
            14'h2805: oData <= 16'h0000;
            14'h2806: oData <= 16'h0000;
            14'h2807: oData <= 16'h0000;
            14'h2808: oData <= 16'h0000;
            14'h2809: oData <= 16'h0000;
            14'h280a: oData <= 16'h0000;
            14'h280b: oData <= 16'h0000;
            14'h280c: oData <= 16'h0000;
            14'h280d: oData <= 16'h0000;
            14'h280e: oData <= 16'h0000;
            14'h280f: oData <= 16'h0000;
            14'h2810: oData <= 16'h0000;
            14'h2811: oData <= 16'h0000;
            14'h2812: oData <= 16'h0000;
            14'h2813: oData <= 16'h0000;
            14'h2814: oData <= 16'h0000;
            14'h2815: oData <= 16'h0000;
            14'h2816: oData <= 16'h0000;
            14'h2817: oData <= 16'h0000;
            14'h2818: oData <= 16'h0000;
            14'h2819: oData <= 16'h0000;
            14'h281a: oData <= 16'h0000;
            14'h281b: oData <= 16'h0000;
            14'h281c: oData <= 16'h0000;
            14'h281d: oData <= 16'h0000;
            14'h281e: oData <= 16'h0000;
            14'h281f: oData <= 16'h0000;
            14'h2820: oData <= 16'h0000;
            14'h2821: oData <= 16'h0000;
            14'h2822: oData <= 16'h0000;
            14'h2823: oData <= 16'h0000;
            14'h2824: oData <= 16'h0000;
            14'h2825: oData <= 16'h0000;
            14'h2826: oData <= 16'h0000;
            14'h2827: oData <= 16'h0000;
            14'h2828: oData <= 16'h0000;
            14'h2829: oData <= 16'h0000;
            14'h282a: oData <= 16'h0000;
            14'h282b: oData <= 16'h0000;
            14'h282c: oData <= 16'h0000;
            14'h282d: oData <= 16'h0000;
            14'h282e: oData <= 16'h0000;
            14'h282f: oData <= 16'h0000;
            14'h2830: oData <= 16'h0000;
            14'h2831: oData <= 16'h0000;
            14'h2832: oData <= 16'h0000;
            14'h2833: oData <= 16'h0000;
            14'h2834: oData <= 16'h0000;
            14'h2835: oData <= 16'h0000;
            14'h2836: oData <= 16'h0000;
            14'h2837: oData <= 16'h0000;
            14'h2838: oData <= 16'h0000;
            14'h2839: oData <= 16'h0000;
            14'h283a: oData <= 16'h0000;
            14'h283b: oData <= 16'h0000;
            14'h283c: oData <= 16'h0000;
            14'h283d: oData <= 16'h0000;
            14'h283e: oData <= 16'h0000;
            14'h283f: oData <= 16'h0000;
            14'h2840: oData <= 16'h0000;
            14'h2841: oData <= 16'h0000;
            14'h2842: oData <= 16'h0000;
            14'h2843: oData <= 16'h0000;
            14'h2844: oData <= 16'h0000;
            14'h2845: oData <= 16'h0000;
            14'h2846: oData <= 16'h0000;
            14'h2847: oData <= 16'h0000;
            14'h2848: oData <= 16'h0000;
            14'h2849: oData <= 16'h0000;
            14'h284a: oData <= 16'h0000;
            14'h284b: oData <= 16'h0000;
            14'h284c: oData <= 16'h0000;
            14'h284d: oData <= 16'h0000;
            14'h284e: oData <= 16'h0000;
            14'h284f: oData <= 16'h0000;
            14'h2850: oData <= 16'h0000;
            14'h2851: oData <= 16'h0000;
            14'h2852: oData <= 16'h0000;
            14'h2853: oData <= 16'h0000;
            14'h2854: oData <= 16'h0000;
            14'h2855: oData <= 16'h0000;
            14'h2856: oData <= 16'h0000;
            14'h2857: oData <= 16'h0000;
            14'h2858: oData <= 16'h0000;
            14'h2859: oData <= 16'h0000;
            14'h285a: oData <= 16'h0000;
            14'h285b: oData <= 16'h0000;
            14'h285c: oData <= 16'h0000;
            14'h285d: oData <= 16'h0000;
            14'h285e: oData <= 16'h0000;
            14'h285f: oData <= 16'h0000;
            14'h2860: oData <= 16'h0000;
            14'h2861: oData <= 16'h0000;
            14'h2862: oData <= 16'h0000;
            14'h2863: oData <= 16'h0000;
            14'h2864: oData <= 16'h0000;
            14'h2865: oData <= 16'h0000;
            14'h2866: oData <= 16'h0000;
            14'h2867: oData <= 16'h0000;
            14'h2868: oData <= 16'h0000;
            14'h2869: oData <= 16'h0000;
            14'h286a: oData <= 16'h0000;
            14'h286b: oData <= 16'h0000;
            14'h286c: oData <= 16'h0000;
            14'h286d: oData <= 16'h0000;
            14'h286e: oData <= 16'h0000;
            14'h286f: oData <= 16'h0000;
            14'h2870: oData <= 16'h0000;
            14'h2871: oData <= 16'h0000;
            14'h2872: oData <= 16'h0000;
            14'h2873: oData <= 16'h0000;
            14'h2874: oData <= 16'h0000;
            14'h2875: oData <= 16'h0000;
            14'h2876: oData <= 16'h0000;
            14'h2877: oData <= 16'h0000;
            14'h2878: oData <= 16'h0000;
            14'h2879: oData <= 16'h0000;
            14'h287a: oData <= 16'h0000;
            14'h287b: oData <= 16'h0000;
            14'h287c: oData <= 16'h0000;
            14'h287d: oData <= 16'h0000;
            14'h287e: oData <= 16'h0000;
            14'h287f: oData <= 16'h0000;
            14'h2880: oData <= 16'h0000;
            14'h2881: oData <= 16'h0000;
            14'h2882: oData <= 16'h0000;
            14'h2883: oData <= 16'h0000;
            14'h2884: oData <= 16'h0000;
            14'h2885: oData <= 16'h0000;
            14'h2886: oData <= 16'h0000;
            14'h2887: oData <= 16'h0000;
            14'h2888: oData <= 16'h0000;
            14'h2889: oData <= 16'h0000;
            14'h288a: oData <= 16'h0000;
            14'h288b: oData <= 16'h0000;
            14'h288c: oData <= 16'h0000;
            14'h288d: oData <= 16'h0000;
            14'h288e: oData <= 16'h0000;
            14'h288f: oData <= 16'h0000;
            14'h2890: oData <= 16'h0000;
            14'h2891: oData <= 16'h0000;
            14'h2892: oData <= 16'h0000;
            14'h2893: oData <= 16'h0000;
            14'h2894: oData <= 16'h0000;
            14'h2895: oData <= 16'h0000;
            14'h2896: oData <= 16'h0000;
            14'h2897: oData <= 16'h0000;
            14'h2898: oData <= 16'h0000;
            14'h2899: oData <= 16'h0000;
            14'h289a: oData <= 16'h0000;
            14'h289b: oData <= 16'h0000;
            14'h289c: oData <= 16'h0000;
            14'h289d: oData <= 16'h0000;
            14'h289e: oData <= 16'h0000;
            14'h289f: oData <= 16'h0000;
            14'h28a0: oData <= 16'h0000;
            14'h28a1: oData <= 16'h0000;
            14'h28a2: oData <= 16'h0000;
            14'h28a3: oData <= 16'h0000;
            14'h28a4: oData <= 16'h0000;
            14'h28a5: oData <= 16'h0000;
            14'h28a6: oData <= 16'h0000;
            14'h28a7: oData <= 16'h0000;
            14'h28a8: oData <= 16'h0000;
            14'h28a9: oData <= 16'h0000;
            14'h28aa: oData <= 16'h0000;
            14'h28ab: oData <= 16'h0000;
            14'h28ac: oData <= 16'h0000;
            14'h28ad: oData <= 16'h0000;
            14'h28ae: oData <= 16'h0000;
            14'h28af: oData <= 16'h0000;
            14'h28b0: oData <= 16'h0000;
            14'h28b1: oData <= 16'h0000;
            14'h28b2: oData <= 16'h0000;
            14'h28b3: oData <= 16'h0000;
            14'h28b4: oData <= 16'h0000;
            14'h28b5: oData <= 16'h0000;
            14'h28b6: oData <= 16'h0000;
            14'h28b7: oData <= 16'h0000;
            14'h28b8: oData <= 16'h0000;
            14'h28b9: oData <= 16'h0000;
            14'h28ba: oData <= 16'h0000;
            14'h28bb: oData <= 16'h0000;
            14'h28bc: oData <= 16'h0000;
            14'h28bd: oData <= 16'h0000;
            14'h28be: oData <= 16'h0000;
            14'h28bf: oData <= 16'h0000;
            14'h28c0: oData <= 16'h0000;
            14'h28c1: oData <= 16'h0000;
            14'h28c2: oData <= 16'h0000;
            14'h28c3: oData <= 16'h0000;
            14'h28c4: oData <= 16'h0000;
            14'h28c5: oData <= 16'h0000;
            14'h28c6: oData <= 16'h0000;
            14'h28c7: oData <= 16'h0000;
            14'h28c8: oData <= 16'h0000;
            14'h28c9: oData <= 16'h0000;
            14'h28ca: oData <= 16'h0000;
            14'h28cb: oData <= 16'h0000;
            14'h28cc: oData <= 16'h0000;
            14'h28cd: oData <= 16'h0000;
            14'h28ce: oData <= 16'h0000;
            14'h28cf: oData <= 16'h0000;
            14'h28d0: oData <= 16'h0000;
            14'h28d1: oData <= 16'h0000;
            14'h28d2: oData <= 16'h0000;
            14'h28d3: oData <= 16'h0000;
            14'h28d4: oData <= 16'h0000;
            14'h28d5: oData <= 16'h0000;
            14'h28d6: oData <= 16'h0000;
            14'h28d7: oData <= 16'h0000;
            14'h28d8: oData <= 16'h0000;
            14'h28d9: oData <= 16'h0000;
            14'h28da: oData <= 16'h0000;
            14'h28db: oData <= 16'h0000;
            14'h28dc: oData <= 16'h0000;
            14'h28dd: oData <= 16'h0000;
            14'h28de: oData <= 16'h0000;
            14'h28df: oData <= 16'h0000;
            14'h28e0: oData <= 16'h0000;
            14'h28e1: oData <= 16'h0000;
            14'h28e2: oData <= 16'h0000;
            14'h28e3: oData <= 16'h0000;
            14'h28e4: oData <= 16'h0000;
            14'h28e5: oData <= 16'h0000;
            14'h28e6: oData <= 16'h0000;
            14'h28e7: oData <= 16'h0000;
            14'h28e8: oData <= 16'h0000;
            14'h28e9: oData <= 16'h0000;
            14'h28ea: oData <= 16'h0000;
            14'h28eb: oData <= 16'h0000;
            14'h28ec: oData <= 16'h0000;
            14'h28ed: oData <= 16'h0000;
            14'h28ee: oData <= 16'h0000;
            14'h28ef: oData <= 16'h0000;
            14'h28f0: oData <= 16'h0000;
            14'h28f1: oData <= 16'h0000;
            14'h28f2: oData <= 16'h0000;
            14'h28f3: oData <= 16'h0000;
            14'h28f4: oData <= 16'h0000;
            14'h28f5: oData <= 16'h0000;
            14'h28f6: oData <= 16'h0000;
            14'h28f7: oData <= 16'h0000;
            14'h28f8: oData <= 16'h0000;
            14'h28f9: oData <= 16'h0000;
            14'h28fa: oData <= 16'h0000;
            14'h28fb: oData <= 16'h0000;
            14'h28fc: oData <= 16'h0000;
            14'h28fd: oData <= 16'h0000;
            14'h28fe: oData <= 16'h0000;
            14'h28ff: oData <= 16'h0000;
            14'h2900: oData <= 16'h0000;
            14'h2901: oData <= 16'h0000;
            14'h2902: oData <= 16'h0000;
            14'h2903: oData <= 16'h0000;
            14'h2904: oData <= 16'h0000;
            14'h2905: oData <= 16'h0000;
            14'h2906: oData <= 16'h0000;
            14'h2907: oData <= 16'h0000;
            14'h2908: oData <= 16'h0000;
            14'h2909: oData <= 16'h0000;
            14'h290a: oData <= 16'h0000;
            14'h290b: oData <= 16'h0000;
            14'h290c: oData <= 16'h0000;
            14'h290d: oData <= 16'h0000;
            14'h290e: oData <= 16'h0000;
            14'h290f: oData <= 16'h0000;
            14'h2910: oData <= 16'h0000;
            14'h2911: oData <= 16'h0000;
            14'h2912: oData <= 16'h0000;
            14'h2913: oData <= 16'h0000;
            14'h2914: oData <= 16'h0000;
            14'h2915: oData <= 16'h0000;
            14'h2916: oData <= 16'h0000;
            14'h2917: oData <= 16'h0000;
            14'h2918: oData <= 16'h0000;
            14'h2919: oData <= 16'h0000;
            14'h291a: oData <= 16'h0000;
            14'h291b: oData <= 16'h0000;
            14'h291c: oData <= 16'h0000;
            14'h291d: oData <= 16'h0000;
            14'h291e: oData <= 16'h0000;
            14'h291f: oData <= 16'h0000;
            14'h2920: oData <= 16'h0000;
            14'h2921: oData <= 16'h0000;
            14'h2922: oData <= 16'h0000;
            14'h2923: oData <= 16'h0000;
            14'h2924: oData <= 16'h0000;
            14'h2925: oData <= 16'h0000;
            14'h2926: oData <= 16'h0000;
            14'h2927: oData <= 16'h0000;
            14'h2928: oData <= 16'h0000;
            14'h2929: oData <= 16'h0000;
            14'h292a: oData <= 16'h0000;
            14'h292b: oData <= 16'h0000;
            14'h292c: oData <= 16'h0000;
            14'h292d: oData <= 16'h0000;
            14'h292e: oData <= 16'h0000;
            14'h292f: oData <= 16'h0000;
            14'h2930: oData <= 16'h0000;
            14'h2931: oData <= 16'h0000;
            14'h2932: oData <= 16'h0000;
            14'h2933: oData <= 16'h0000;
            14'h2934: oData <= 16'h0000;
            14'h2935: oData <= 16'h0000;
            14'h2936: oData <= 16'h0000;
            14'h2937: oData <= 16'h0000;
            14'h2938: oData <= 16'h0000;
            14'h2939: oData <= 16'h0000;
            14'h293a: oData <= 16'h0000;
            14'h293b: oData <= 16'h0000;
            14'h293c: oData <= 16'h0000;
            14'h293d: oData <= 16'h0000;
            14'h293e: oData <= 16'h0000;
            14'h293f: oData <= 16'h0000;
            14'h2940: oData <= 16'h0000;
            14'h2941: oData <= 16'h0000;
            14'h2942: oData <= 16'h0000;
            14'h2943: oData <= 16'h0000;
            14'h2944: oData <= 16'h0000;
            14'h2945: oData <= 16'h0000;
            14'h2946: oData <= 16'h0000;
            14'h2947: oData <= 16'h0000;
            14'h2948: oData <= 16'h0000;
            14'h2949: oData <= 16'h0000;
            14'h294a: oData <= 16'h0000;
            14'h294b: oData <= 16'h0000;
            14'h294c: oData <= 16'h0000;
            14'h294d: oData <= 16'h0000;
            14'h294e: oData <= 16'h0000;
            14'h294f: oData <= 16'h0000;
            14'h2950: oData <= 16'h0000;
            14'h2951: oData <= 16'h0000;
            14'h2952: oData <= 16'h0000;
            14'h2953: oData <= 16'h0000;
            14'h2954: oData <= 16'h0000;
            14'h2955: oData <= 16'h0000;
            14'h2956: oData <= 16'h0000;
            14'h2957: oData <= 16'h0000;
            14'h2958: oData <= 16'h0000;
            14'h2959: oData <= 16'h0000;
            14'h295a: oData <= 16'h0000;
            14'h295b: oData <= 16'h0000;
            14'h295c: oData <= 16'h0000;
            14'h295d: oData <= 16'h0000;
            14'h295e: oData <= 16'h0000;
            14'h295f: oData <= 16'h0000;
            14'h2960: oData <= 16'h0000;
            14'h2961: oData <= 16'h0000;
            14'h2962: oData <= 16'h0000;
            14'h2963: oData <= 16'h0000;
            14'h2964: oData <= 16'h0000;
            14'h2965: oData <= 16'h0000;
            14'h2966: oData <= 16'h0000;
            14'h2967: oData <= 16'h0000;
            14'h2968: oData <= 16'h0000;
            14'h2969: oData <= 16'h0000;
            14'h296a: oData <= 16'h0000;
            14'h296b: oData <= 16'h0000;
            14'h296c: oData <= 16'h0000;
            14'h296d: oData <= 16'h0000;
            14'h296e: oData <= 16'h0000;
            14'h296f: oData <= 16'h0000;
            14'h2970: oData <= 16'h0000;
            14'h2971: oData <= 16'h0000;
            14'h2972: oData <= 16'h0000;
            14'h2973: oData <= 16'h0000;
            14'h2974: oData <= 16'h0000;
            14'h2975: oData <= 16'h0000;
            14'h2976: oData <= 16'h0000;
            14'h2977: oData <= 16'h0000;
            14'h2978: oData <= 16'h0000;
            14'h2979: oData <= 16'h0000;
            14'h297a: oData <= 16'h0000;
            14'h297b: oData <= 16'h0000;
            14'h297c: oData <= 16'h0000;
            14'h297d: oData <= 16'h0000;
            14'h297e: oData <= 16'h0000;
            14'h297f: oData <= 16'h0000;
            14'h2980: oData <= 16'h0000;
            14'h2981: oData <= 16'h0000;
            14'h2982: oData <= 16'h0000;
            14'h2983: oData <= 16'h0000;
            14'h2984: oData <= 16'h0000;
            14'h2985: oData <= 16'h0000;
            14'h2986: oData <= 16'h0000;
            14'h2987: oData <= 16'h0000;
            14'h2988: oData <= 16'h0000;
            14'h2989: oData <= 16'h0000;
            14'h298a: oData <= 16'h0000;
            14'h298b: oData <= 16'h0000;
            14'h298c: oData <= 16'h0000;
            14'h298d: oData <= 16'h0000;
            14'h298e: oData <= 16'h0000;
            14'h298f: oData <= 16'h0000;
            14'h2990: oData <= 16'h0000;
            14'h2991: oData <= 16'h0000;
            14'h2992: oData <= 16'h0000;
            14'h2993: oData <= 16'h0000;
            14'h2994: oData <= 16'h0000;
            14'h2995: oData <= 16'h0000;
            14'h2996: oData <= 16'h0000;
            14'h2997: oData <= 16'h0000;
            14'h2998: oData <= 16'h0000;
            14'h2999: oData <= 16'h0000;
            14'h299a: oData <= 16'h0000;
            14'h299b: oData <= 16'h0000;
            14'h299c: oData <= 16'h0000;
            14'h299d: oData <= 16'h0000;
            14'h299e: oData <= 16'h0000;
            14'h299f: oData <= 16'h0000;
            14'h29a0: oData <= 16'h0000;
            14'h29a1: oData <= 16'h0000;
            14'h29a2: oData <= 16'h0000;
            14'h29a3: oData <= 16'h0000;
            14'h29a4: oData <= 16'h0000;
            14'h29a5: oData <= 16'h0000;
            14'h29a6: oData <= 16'h0000;
            14'h29a7: oData <= 16'h0000;
            14'h29a8: oData <= 16'h0000;
            14'h29a9: oData <= 16'h0000;
            14'h29aa: oData <= 16'h0000;
            14'h29ab: oData <= 16'h0000;
            14'h29ac: oData <= 16'h0000;
            14'h29ad: oData <= 16'h0000;
            14'h29ae: oData <= 16'h0000;
            14'h29af: oData <= 16'h0000;
            14'h29b0: oData <= 16'h0000;
            14'h29b1: oData <= 16'h0000;
            14'h29b2: oData <= 16'h0000;
            14'h29b3: oData <= 16'h0000;
            14'h29b4: oData <= 16'h0000;
            14'h29b5: oData <= 16'h0000;
            14'h29b6: oData <= 16'h0000;
            14'h29b7: oData <= 16'h0000;
            14'h29b8: oData <= 16'h0000;
            14'h29b9: oData <= 16'h0000;
            14'h29ba: oData <= 16'h0000;
            14'h29bb: oData <= 16'h0000;
            14'h29bc: oData <= 16'h0000;
            14'h29bd: oData <= 16'h0000;
            14'h29be: oData <= 16'h0000;
            14'h29bf: oData <= 16'h0000;
            14'h29c0: oData <= 16'h0000;
            14'h29c1: oData <= 16'h0000;
            14'h29c2: oData <= 16'h0000;
            14'h29c3: oData <= 16'h0000;
            14'h29c4: oData <= 16'h0000;
            14'h29c5: oData <= 16'h0000;
            14'h29c6: oData <= 16'h0000;
            14'h29c7: oData <= 16'h0000;
            14'h29c8: oData <= 16'h0000;
            14'h29c9: oData <= 16'h0000;
            14'h29ca: oData <= 16'h0000;
            14'h29cb: oData <= 16'h0000;
            14'h29cc: oData <= 16'h0000;
            14'h29cd: oData <= 16'h0000;
            14'h29ce: oData <= 16'h0000;
            14'h29cf: oData <= 16'h0000;
            14'h29d0: oData <= 16'h0000;
            14'h29d1: oData <= 16'h0000;
            14'h29d2: oData <= 16'h0000;
            14'h29d3: oData <= 16'h0000;
            14'h29d4: oData <= 16'h0000;
            14'h29d5: oData <= 16'h0000;
            14'h29d6: oData <= 16'h0000;
            14'h29d7: oData <= 16'h0000;
            14'h29d8: oData <= 16'h0000;
            14'h29d9: oData <= 16'h0000;
            14'h29da: oData <= 16'h0000;
            14'h29db: oData <= 16'h0000;
            14'h29dc: oData <= 16'h0000;
            14'h29dd: oData <= 16'h0000;
            14'h29de: oData <= 16'h0000;
            14'h29df: oData <= 16'h0000;
            14'h29e0: oData <= 16'h0000;
            14'h29e1: oData <= 16'h0000;
            14'h29e2: oData <= 16'h0000;
            14'h29e3: oData <= 16'h0000;
            14'h29e4: oData <= 16'h0000;
            14'h29e5: oData <= 16'h0000;
            14'h29e6: oData <= 16'h0000;
            14'h29e7: oData <= 16'h0000;
            14'h29e8: oData <= 16'h0000;
            14'h29e9: oData <= 16'h0000;
            14'h29ea: oData <= 16'h0000;
            14'h29eb: oData <= 16'h0000;
            14'h29ec: oData <= 16'h0000;
            14'h29ed: oData <= 16'h0000;
            14'h29ee: oData <= 16'h0000;
            14'h29ef: oData <= 16'h0000;
            14'h29f0: oData <= 16'h0000;
            14'h29f1: oData <= 16'h0000;
            14'h29f2: oData <= 16'h0000;
            14'h29f3: oData <= 16'h0000;
            14'h29f4: oData <= 16'h0000;
            14'h29f5: oData <= 16'h0000;
            14'h29f6: oData <= 16'h0000;
            14'h29f7: oData <= 16'h0000;
            14'h29f8: oData <= 16'h0000;
            14'h29f9: oData <= 16'h0000;
            14'h29fa: oData <= 16'h0000;
            14'h29fb: oData <= 16'h0000;
            14'h29fc: oData <= 16'h0000;
            14'h29fd: oData <= 16'h0000;
            14'h29fe: oData <= 16'h0000;
            14'h29ff: oData <= 16'h0000;
            14'h2a00: oData <= 16'h0000;
            14'h2a01: oData <= 16'h0000;
            14'h2a02: oData <= 16'h0000;
            14'h2a03: oData <= 16'h0000;
            14'h2a04: oData <= 16'h0000;
            14'h2a05: oData <= 16'h0000;
            14'h2a06: oData <= 16'h0000;
            14'h2a07: oData <= 16'h0000;
            14'h2a08: oData <= 16'h0000;
            14'h2a09: oData <= 16'h0000;
            14'h2a0a: oData <= 16'h0000;
            14'h2a0b: oData <= 16'h0000;
            14'h2a0c: oData <= 16'h0000;
            14'h2a0d: oData <= 16'h0000;
            14'h2a0e: oData <= 16'h0000;
            14'h2a0f: oData <= 16'h0000;
            14'h2a10: oData <= 16'h0000;
            14'h2a11: oData <= 16'h0000;
            14'h2a12: oData <= 16'h0000;
            14'h2a13: oData <= 16'h0000;
            14'h2a14: oData <= 16'h0000;
            14'h2a15: oData <= 16'h0000;
            14'h2a16: oData <= 16'h0000;
            14'h2a17: oData <= 16'h0000;
            14'h2a18: oData <= 16'h0000;
            14'h2a19: oData <= 16'h0000;
            14'h2a1a: oData <= 16'h0000;
            14'h2a1b: oData <= 16'h0000;
            14'h2a1c: oData <= 16'h0000;
            14'h2a1d: oData <= 16'h0000;
            14'h2a1e: oData <= 16'h0000;
            14'h2a1f: oData <= 16'h0000;
            14'h2a20: oData <= 16'h0000;
            14'h2a21: oData <= 16'h0000;
            14'h2a22: oData <= 16'h0000;
            14'h2a23: oData <= 16'h0000;
            14'h2a24: oData <= 16'h0000;
            14'h2a25: oData <= 16'h0000;
            14'h2a26: oData <= 16'h0000;
            14'h2a27: oData <= 16'h0000;
            14'h2a28: oData <= 16'h0000;
            14'h2a29: oData <= 16'h0000;
            14'h2a2a: oData <= 16'h0000;
            14'h2a2b: oData <= 16'h0000;
            14'h2a2c: oData <= 16'h0000;
            14'h2a2d: oData <= 16'h0000;
            14'h2a2e: oData <= 16'h0000;
            14'h2a2f: oData <= 16'h0000;
            14'h2a30: oData <= 16'h0000;
            14'h2a31: oData <= 16'h0000;
            14'h2a32: oData <= 16'h0000;
            14'h2a33: oData <= 16'h0000;
            14'h2a34: oData <= 16'h0000;
            14'h2a35: oData <= 16'h0000;
            14'h2a36: oData <= 16'h0000;
            14'h2a37: oData <= 16'h0000;
            14'h2a38: oData <= 16'h0000;
            14'h2a39: oData <= 16'h0000;
            14'h2a3a: oData <= 16'h0000;
            14'h2a3b: oData <= 16'h0000;
            14'h2a3c: oData <= 16'h0000;
            14'h2a3d: oData <= 16'h0000;
            14'h2a3e: oData <= 16'h0000;
            14'h2a3f: oData <= 16'h0000;
            14'h2a40: oData <= 16'h0000;
            14'h2a41: oData <= 16'h0000;
            14'h2a42: oData <= 16'h0000;
            14'h2a43: oData <= 16'h0000;
            14'h2a44: oData <= 16'h0000;
            14'h2a45: oData <= 16'h0000;
            14'h2a46: oData <= 16'h0000;
            14'h2a47: oData <= 16'h0000;
            14'h2a48: oData <= 16'h0000;
            14'h2a49: oData <= 16'h0000;
            14'h2a4a: oData <= 16'h0000;
            14'h2a4b: oData <= 16'h0000;
            14'h2a4c: oData <= 16'h0000;
            14'h2a4d: oData <= 16'h0000;
            14'h2a4e: oData <= 16'h0000;
            14'h2a4f: oData <= 16'h0000;
            14'h2a50: oData <= 16'h0000;
            14'h2a51: oData <= 16'h0000;
            14'h2a52: oData <= 16'h0000;
            14'h2a53: oData <= 16'h0000;
            14'h2a54: oData <= 16'h0000;
            14'h2a55: oData <= 16'h0000;
            14'h2a56: oData <= 16'h0000;
            14'h2a57: oData <= 16'h0000;
            14'h2a58: oData <= 16'h0000;
            14'h2a59: oData <= 16'h0000;
            14'h2a5a: oData <= 16'h0000;
            14'h2a5b: oData <= 16'h0000;
            14'h2a5c: oData <= 16'h0000;
            14'h2a5d: oData <= 16'h0000;
            14'h2a5e: oData <= 16'h0000;
            14'h2a5f: oData <= 16'h0000;
            14'h2a60: oData <= 16'h0000;
            14'h2a61: oData <= 16'h0000;
            14'h2a62: oData <= 16'h0000;
            14'h2a63: oData <= 16'h0000;
            14'h2a64: oData <= 16'h0000;
            14'h2a65: oData <= 16'h0000;
            14'h2a66: oData <= 16'h0000;
            14'h2a67: oData <= 16'h0000;
            14'h2a68: oData <= 16'h0000;
            14'h2a69: oData <= 16'h0000;
            14'h2a6a: oData <= 16'h0000;
            14'h2a6b: oData <= 16'h0000;
            14'h2a6c: oData <= 16'h0000;
            14'h2a6d: oData <= 16'h0000;
            14'h2a6e: oData <= 16'h0000;
            14'h2a6f: oData <= 16'h0000;
            14'h2a70: oData <= 16'h0000;
            14'h2a71: oData <= 16'h0000;
            14'h2a72: oData <= 16'h0000;
            14'h2a73: oData <= 16'h0000;
            14'h2a74: oData <= 16'h0000;
            14'h2a75: oData <= 16'h0000;
            14'h2a76: oData <= 16'h0000;
            14'h2a77: oData <= 16'h0000;
            14'h2a78: oData <= 16'h0000;
            14'h2a79: oData <= 16'h0000;
            14'h2a7a: oData <= 16'h0000;
            14'h2a7b: oData <= 16'h0000;
            14'h2a7c: oData <= 16'h0000;
            14'h2a7d: oData <= 16'h0000;
            14'h2a7e: oData <= 16'h0000;
            14'h2a7f: oData <= 16'h0000;
            14'h2a80: oData <= 16'h0000;
            14'h2a81: oData <= 16'h0000;
            14'h2a82: oData <= 16'h0000;
            14'h2a83: oData <= 16'h0000;
            14'h2a84: oData <= 16'h0000;
            14'h2a85: oData <= 16'h0000;
            14'h2a86: oData <= 16'h0000;
            14'h2a87: oData <= 16'h0000;
            14'h2a88: oData <= 16'h0000;
            14'h2a89: oData <= 16'h0000;
            14'h2a8a: oData <= 16'h0000;
            14'h2a8b: oData <= 16'h0000;
            14'h2a8c: oData <= 16'h0000;
            14'h2a8d: oData <= 16'h0000;
            14'h2a8e: oData <= 16'h0000;
            14'h2a8f: oData <= 16'h0000;
            14'h2a90: oData <= 16'h0000;
            14'h2a91: oData <= 16'h0000;
            14'h2a92: oData <= 16'h0000;
            14'h2a93: oData <= 16'h0000;
            14'h2a94: oData <= 16'h0000;
            14'h2a95: oData <= 16'h0000;
            14'h2a96: oData <= 16'h0000;
            14'h2a97: oData <= 16'h0000;
            14'h2a98: oData <= 16'h0000;
            14'h2a99: oData <= 16'h0000;
            14'h2a9a: oData <= 16'h0000;
            14'h2a9b: oData <= 16'h0000;
            14'h2a9c: oData <= 16'h0000;
            14'h2a9d: oData <= 16'h0000;
            14'h2a9e: oData <= 16'h0000;
            14'h2a9f: oData <= 16'h0000;
            14'h2aa0: oData <= 16'h0000;
            14'h2aa1: oData <= 16'h0000;
            14'h2aa2: oData <= 16'h0000;
            14'h2aa3: oData <= 16'h0000;
            14'h2aa4: oData <= 16'h0000;
            14'h2aa5: oData <= 16'h0000;
            14'h2aa6: oData <= 16'h0000;
            14'h2aa7: oData <= 16'h0000;
            14'h2aa8: oData <= 16'h0000;
            14'h2aa9: oData <= 16'h0000;
            14'h2aaa: oData <= 16'h0000;
            14'h2aab: oData <= 16'h0000;
            14'h2aac: oData <= 16'h0000;
            14'h2aad: oData <= 16'h0000;
            14'h2aae: oData <= 16'h0000;
            14'h2aaf: oData <= 16'h0000;
            14'h2ab0: oData <= 16'h0000;
            14'h2ab1: oData <= 16'h0000;
            14'h2ab2: oData <= 16'h0000;
            14'h2ab3: oData <= 16'h0000;
            14'h2ab4: oData <= 16'h0000;
            14'h2ab5: oData <= 16'h0000;
            14'h2ab6: oData <= 16'h0000;
            14'h2ab7: oData <= 16'h0000;
            14'h2ab8: oData <= 16'h0000;
            14'h2ab9: oData <= 16'h0000;
            14'h2aba: oData <= 16'h0000;
            14'h2abb: oData <= 16'h0000;
            14'h2abc: oData <= 16'h0000;
            14'h2abd: oData <= 16'h0000;
            14'h2abe: oData <= 16'h0000;
            14'h2abf: oData <= 16'h0000;
            14'h2ac0: oData <= 16'h0000;
            14'h2ac1: oData <= 16'h0000;
            14'h2ac2: oData <= 16'h0000;
            14'h2ac3: oData <= 16'h0000;
            14'h2ac4: oData <= 16'h0000;
            14'h2ac5: oData <= 16'h0000;
            14'h2ac6: oData <= 16'h0000;
            14'h2ac7: oData <= 16'h0000;
            14'h2ac8: oData <= 16'h0000;
            14'h2ac9: oData <= 16'h0000;
            14'h2aca: oData <= 16'h0000;
            14'h2acb: oData <= 16'h0000;
            14'h2acc: oData <= 16'h0000;
            14'h2acd: oData <= 16'h0000;
            14'h2ace: oData <= 16'h0000;
            14'h2acf: oData <= 16'h0000;
            14'h2ad0: oData <= 16'h0000;
            14'h2ad1: oData <= 16'h0000;
            14'h2ad2: oData <= 16'h0000;
            14'h2ad3: oData <= 16'h0000;
            14'h2ad4: oData <= 16'h0000;
            14'h2ad5: oData <= 16'h0000;
            14'h2ad6: oData <= 16'h0000;
            14'h2ad7: oData <= 16'h0000;
            14'h2ad8: oData <= 16'h0000;
            14'h2ad9: oData <= 16'h0000;
            14'h2ada: oData <= 16'h0000;
            14'h2adb: oData <= 16'h0000;
            14'h2adc: oData <= 16'h0000;
            14'h2add: oData <= 16'h0000;
            14'h2ade: oData <= 16'h0000;
            14'h2adf: oData <= 16'h0000;
            14'h2ae0: oData <= 16'h0000;
            14'h2ae1: oData <= 16'h0000;
            14'h2ae2: oData <= 16'h0000;
            14'h2ae3: oData <= 16'h0000;
            14'h2ae4: oData <= 16'h0000;
            14'h2ae5: oData <= 16'h0000;
            14'h2ae6: oData <= 16'h0000;
            14'h2ae7: oData <= 16'h0000;
            14'h2ae8: oData <= 16'h0000;
            14'h2ae9: oData <= 16'h0000;
            14'h2aea: oData <= 16'h0000;
            14'h2aeb: oData <= 16'h0000;
            14'h2aec: oData <= 16'h0000;
            14'h2aed: oData <= 16'h0000;
            14'h2aee: oData <= 16'h0000;
            14'h2aef: oData <= 16'h0000;
            14'h2af0: oData <= 16'h0000;
            14'h2af1: oData <= 16'h0000;
            14'h2af2: oData <= 16'h0000;
            14'h2af3: oData <= 16'h0000;
            14'h2af4: oData <= 16'h0000;
            14'h2af5: oData <= 16'h0000;
            14'h2af6: oData <= 16'h0000;
            14'h2af7: oData <= 16'h0000;
            14'h2af8: oData <= 16'h0000;
            14'h2af9: oData <= 16'h0000;
            14'h2afa: oData <= 16'h0000;
            14'h2afb: oData <= 16'h0000;
            14'h2afc: oData <= 16'h0000;
            14'h2afd: oData <= 16'h0000;
            14'h2afe: oData <= 16'h0000;
            14'h2aff: oData <= 16'h0000;
            14'h2b00: oData <= 16'h0000;
            14'h2b01: oData <= 16'h0000;
            14'h2b02: oData <= 16'h0000;
            14'h2b03: oData <= 16'h0000;
            14'h2b04: oData <= 16'h0000;
            14'h2b05: oData <= 16'h0000;
            14'h2b06: oData <= 16'h0000;
            14'h2b07: oData <= 16'h0000;
            14'h2b08: oData <= 16'h0000;
            14'h2b09: oData <= 16'h0000;
            14'h2b0a: oData <= 16'h0000;
            14'h2b0b: oData <= 16'h0000;
            14'h2b0c: oData <= 16'h0000;
            14'h2b0d: oData <= 16'h0000;
            14'h2b0e: oData <= 16'h0000;
            14'h2b0f: oData <= 16'h0000;
            14'h2b10: oData <= 16'h0000;
            14'h2b11: oData <= 16'h0000;
            14'h2b12: oData <= 16'h0000;
            14'h2b13: oData <= 16'h0000;
            14'h2b14: oData <= 16'h0000;
            14'h2b15: oData <= 16'h0000;
            14'h2b16: oData <= 16'h0000;
            14'h2b17: oData <= 16'h0000;
            14'h2b18: oData <= 16'h0000;
            14'h2b19: oData <= 16'h0000;
            14'h2b1a: oData <= 16'h0000;
            14'h2b1b: oData <= 16'h0000;
            14'h2b1c: oData <= 16'h0000;
            14'h2b1d: oData <= 16'h0000;
            14'h2b1e: oData <= 16'h0000;
            14'h2b1f: oData <= 16'h0000;
            14'h2b20: oData <= 16'h0000;
            14'h2b21: oData <= 16'h0000;
            14'h2b22: oData <= 16'h0000;
            14'h2b23: oData <= 16'h0000;
            14'h2b24: oData <= 16'h0000;
            14'h2b25: oData <= 16'h0000;
            14'h2b26: oData <= 16'h0000;
            14'h2b27: oData <= 16'h0000;
            14'h2b28: oData <= 16'h0000;
            14'h2b29: oData <= 16'h0000;
            14'h2b2a: oData <= 16'h0000;
            14'h2b2b: oData <= 16'h0000;
            14'h2b2c: oData <= 16'h0000;
            14'h2b2d: oData <= 16'h0000;
            14'h2b2e: oData <= 16'h0000;
            14'h2b2f: oData <= 16'h0000;
            14'h2b30: oData <= 16'h0000;
            14'h2b31: oData <= 16'h0000;
            14'h2b32: oData <= 16'h0000;
            14'h2b33: oData <= 16'h0000;
            14'h2b34: oData <= 16'h0000;
            14'h2b35: oData <= 16'h0000;
            14'h2b36: oData <= 16'h0000;
            14'h2b37: oData <= 16'h0000;
            14'h2b38: oData <= 16'h0000;
            14'h2b39: oData <= 16'h0000;
            14'h2b3a: oData <= 16'h0000;
            14'h2b3b: oData <= 16'h0000;
            14'h2b3c: oData <= 16'h0000;
            14'h2b3d: oData <= 16'h0000;
            14'h2b3e: oData <= 16'h0000;
            14'h2b3f: oData <= 16'h0000;
            14'h2b40: oData <= 16'h0000;
            14'h2b41: oData <= 16'h0000;
            14'h2b42: oData <= 16'h0000;
            14'h2b43: oData <= 16'h0000;
            14'h2b44: oData <= 16'h0000;
            14'h2b45: oData <= 16'h0000;
            14'h2b46: oData <= 16'h0000;
            14'h2b47: oData <= 16'h0000;
            14'h2b48: oData <= 16'h0000;
            14'h2b49: oData <= 16'h0000;
            14'h2b4a: oData <= 16'h0000;
            14'h2b4b: oData <= 16'h0000;
            14'h2b4c: oData <= 16'h0000;
            14'h2b4d: oData <= 16'h0000;
            14'h2b4e: oData <= 16'h0000;
            14'h2b4f: oData <= 16'h0000;
            14'h2b50: oData <= 16'h0000;
            14'h2b51: oData <= 16'h0000;
            14'h2b52: oData <= 16'h0000;
            14'h2b53: oData <= 16'h0000;
            14'h2b54: oData <= 16'h0000;
            14'h2b55: oData <= 16'h0000;
            14'h2b56: oData <= 16'h0000;
            14'h2b57: oData <= 16'h0000;
            14'h2b58: oData <= 16'h0000;
            14'h2b59: oData <= 16'h0000;
            14'h2b5a: oData <= 16'h0000;
            14'h2b5b: oData <= 16'h0000;
            14'h2b5c: oData <= 16'h0000;
            14'h2b5d: oData <= 16'h0000;
            14'h2b5e: oData <= 16'h0000;
            14'h2b5f: oData <= 16'h0000;
            14'h2b60: oData <= 16'h0000;
            14'h2b61: oData <= 16'h0000;
            14'h2b62: oData <= 16'h0000;
            14'h2b63: oData <= 16'h0000;
            14'h2b64: oData <= 16'h0000;
            14'h2b65: oData <= 16'h0000;
            14'h2b66: oData <= 16'h0000;
            14'h2b67: oData <= 16'h0000;
            14'h2b68: oData <= 16'h0000;
            14'h2b69: oData <= 16'h0000;
            14'h2b6a: oData <= 16'h0000;
            14'h2b6b: oData <= 16'h0000;
            14'h2b6c: oData <= 16'h0000;
            14'h2b6d: oData <= 16'h0000;
            14'h2b6e: oData <= 16'h0000;
            14'h2b6f: oData <= 16'h0000;
            14'h2b70: oData <= 16'h0000;
            14'h2b71: oData <= 16'h0000;
            14'h2b72: oData <= 16'h0000;
            14'h2b73: oData <= 16'h0000;
            14'h2b74: oData <= 16'h0000;
            14'h2b75: oData <= 16'h0000;
            14'h2b76: oData <= 16'h0000;
            14'h2b77: oData <= 16'h0000;
            14'h2b78: oData <= 16'h0000;
            14'h2b79: oData <= 16'h0000;
            14'h2b7a: oData <= 16'h0000;
            14'h2b7b: oData <= 16'h0000;
            14'h2b7c: oData <= 16'h0000;
            14'h2b7d: oData <= 16'h0000;
            14'h2b7e: oData <= 16'h0000;
            14'h2b7f: oData <= 16'h0000;
            14'h2b80: oData <= 16'h0000;
            14'h2b81: oData <= 16'h0000;
            14'h2b82: oData <= 16'h0000;
            14'h2b83: oData <= 16'h0000;
            14'h2b84: oData <= 16'h0000;
            14'h2b85: oData <= 16'h0000;
            14'h2b86: oData <= 16'h0000;
            14'h2b87: oData <= 16'h0000;
            14'h2b88: oData <= 16'h0000;
            14'h2b89: oData <= 16'h0000;
            14'h2b8a: oData <= 16'h0000;
            14'h2b8b: oData <= 16'h0000;
            14'h2b8c: oData <= 16'h0000;
            14'h2b8d: oData <= 16'h0000;
            14'h2b8e: oData <= 16'h0000;
            14'h2b8f: oData <= 16'h0000;
            14'h2b90: oData <= 16'h0000;
            14'h2b91: oData <= 16'h0000;
            14'h2b92: oData <= 16'h0000;
            14'h2b93: oData <= 16'h0000;
            14'h2b94: oData <= 16'h0000;
            14'h2b95: oData <= 16'h0000;
            14'h2b96: oData <= 16'h0000;
            14'h2b97: oData <= 16'h0000;
            14'h2b98: oData <= 16'h0000;
            14'h2b99: oData <= 16'h0000;
            14'h2b9a: oData <= 16'h0000;
            14'h2b9b: oData <= 16'h0000;
            14'h2b9c: oData <= 16'h0000;
            14'h2b9d: oData <= 16'h0000;
            14'h2b9e: oData <= 16'h0000;
            14'h2b9f: oData <= 16'h0000;
            14'h2ba0: oData <= 16'h0000;
            14'h2ba1: oData <= 16'h0000;
            14'h2ba2: oData <= 16'h0000;
            14'h2ba3: oData <= 16'h0000;
            14'h2ba4: oData <= 16'h0000;
            14'h2ba5: oData <= 16'h0000;
            14'h2ba6: oData <= 16'h0000;
            14'h2ba7: oData <= 16'h0000;
            14'h2ba8: oData <= 16'h0000;
            14'h2ba9: oData <= 16'h0000;
            14'h2baa: oData <= 16'h0000;
            14'h2bab: oData <= 16'h0000;
            14'h2bac: oData <= 16'h0000;
            14'h2bad: oData <= 16'h0000;
            14'h2bae: oData <= 16'h0000;
            14'h2baf: oData <= 16'h0000;
            14'h2bb0: oData <= 16'h0000;
            14'h2bb1: oData <= 16'h0000;
            14'h2bb2: oData <= 16'h0000;
            14'h2bb3: oData <= 16'h0000;
            14'h2bb4: oData <= 16'h0000;
            14'h2bb5: oData <= 16'h0000;
            14'h2bb6: oData <= 16'h0000;
            14'h2bb7: oData <= 16'h0000;
            14'h2bb8: oData <= 16'h0000;
            14'h2bb9: oData <= 16'h0000;
            14'h2bba: oData <= 16'h0000;
            14'h2bbb: oData <= 16'h0000;
            14'h2bbc: oData <= 16'h0000;
            14'h2bbd: oData <= 16'h0000;
            14'h2bbe: oData <= 16'h0000;
            14'h2bbf: oData <= 16'h0000;
            14'h2bc0: oData <= 16'h0000;
            14'h2bc1: oData <= 16'h0000;
            14'h2bc2: oData <= 16'h0000;
            14'h2bc3: oData <= 16'h0000;
            14'h2bc4: oData <= 16'h0000;
            14'h2bc5: oData <= 16'h0000;
            14'h2bc6: oData <= 16'h0000;
            14'h2bc7: oData <= 16'h0000;
            14'h2bc8: oData <= 16'h0000;
            14'h2bc9: oData <= 16'h0000;
            14'h2bca: oData <= 16'h0000;
            14'h2bcb: oData <= 16'h0000;
            14'h2bcc: oData <= 16'h0000;
            14'h2bcd: oData <= 16'h0000;
            14'h2bce: oData <= 16'h0000;
            14'h2bcf: oData <= 16'h0000;
            14'h2bd0: oData <= 16'h0000;
            14'h2bd1: oData <= 16'h0000;
            14'h2bd2: oData <= 16'h0000;
            14'h2bd3: oData <= 16'h0000;
            14'h2bd4: oData <= 16'h0000;
            14'h2bd5: oData <= 16'h0000;
            14'h2bd6: oData <= 16'h0000;
            14'h2bd7: oData <= 16'h0000;
            14'h2bd8: oData <= 16'h0000;
            14'h2bd9: oData <= 16'h0000;
            14'h2bda: oData <= 16'h0000;
            14'h2bdb: oData <= 16'h0000;
            14'h2bdc: oData <= 16'h0000;
            14'h2bdd: oData <= 16'h0000;
            14'h2bde: oData <= 16'h0000;
            14'h2bdf: oData <= 16'h0000;
            14'h2be0: oData <= 16'h0000;
            14'h2be1: oData <= 16'h0000;
            14'h2be2: oData <= 16'h0000;
            14'h2be3: oData <= 16'h0000;
            14'h2be4: oData <= 16'h0000;
            14'h2be5: oData <= 16'h0000;
            14'h2be6: oData <= 16'h0000;
            14'h2be7: oData <= 16'h0000;
            14'h2be8: oData <= 16'h0000;
            14'h2be9: oData <= 16'h0000;
            14'h2bea: oData <= 16'h0000;
            14'h2beb: oData <= 16'h0000;
            14'h2bec: oData <= 16'h0000;
            14'h2bed: oData <= 16'h0000;
            14'h2bee: oData <= 16'h0000;
            14'h2bef: oData <= 16'h0000;
            14'h2bf0: oData <= 16'h0000;
            14'h2bf1: oData <= 16'h0000;
            14'h2bf2: oData <= 16'h0000;
            14'h2bf3: oData <= 16'h0000;
            14'h2bf4: oData <= 16'h0000;
            14'h2bf5: oData <= 16'h0000;
            14'h2bf6: oData <= 16'h0000;
            14'h2bf7: oData <= 16'h0000;
            14'h2bf8: oData <= 16'h0000;
            14'h2bf9: oData <= 16'h0000;
            14'h2bfa: oData <= 16'h0000;
            14'h2bfb: oData <= 16'h0000;
            14'h2bfc: oData <= 16'h0000;
            14'h2bfd: oData <= 16'h0000;
            14'h2bfe: oData <= 16'h0000;
            14'h2bff: oData <= 16'h0000;
            14'h2c00: oData <= 16'h0000;
            14'h2c01: oData <= 16'h0000;
            14'h2c02: oData <= 16'h0000;
            14'h2c03: oData <= 16'h0000;
            14'h2c04: oData <= 16'h0000;
            14'h2c05: oData <= 16'h0000;
            14'h2c06: oData <= 16'h0000;
            14'h2c07: oData <= 16'h0000;
            14'h2c08: oData <= 16'h0000;
            14'h2c09: oData <= 16'h0000;
            14'h2c0a: oData <= 16'h0000;
            14'h2c0b: oData <= 16'h0000;
            14'h2c0c: oData <= 16'h0000;
            14'h2c0d: oData <= 16'h0000;
            14'h2c0e: oData <= 16'h0000;
            14'h2c0f: oData <= 16'h0000;
            14'h2c10: oData <= 16'h0000;
            14'h2c11: oData <= 16'h0000;
            14'h2c12: oData <= 16'h0000;
            14'h2c13: oData <= 16'h0000;
            14'h2c14: oData <= 16'h0000;
            14'h2c15: oData <= 16'h0000;
            14'h2c16: oData <= 16'h0000;
            14'h2c17: oData <= 16'h0000;
            14'h2c18: oData <= 16'h0000;
            14'h2c19: oData <= 16'h0000;
            14'h2c1a: oData <= 16'h0000;
            14'h2c1b: oData <= 16'h0000;
            14'h2c1c: oData <= 16'h0000;
            14'h2c1d: oData <= 16'h0000;
            14'h2c1e: oData <= 16'h0000;
            14'h2c1f: oData <= 16'h0000;
            14'h2c20: oData <= 16'h0000;
            14'h2c21: oData <= 16'h0000;
            14'h2c22: oData <= 16'h0000;
            14'h2c23: oData <= 16'h0000;
            14'h2c24: oData <= 16'h0000;
            14'h2c25: oData <= 16'h0000;
            14'h2c26: oData <= 16'h0000;
            14'h2c27: oData <= 16'h0000;
            14'h2c28: oData <= 16'h0000;
            14'h2c29: oData <= 16'h0000;
            14'h2c2a: oData <= 16'h0000;
            14'h2c2b: oData <= 16'h0000;
            14'h2c2c: oData <= 16'h0000;
            14'h2c2d: oData <= 16'h0000;
            14'h2c2e: oData <= 16'h0000;
            14'h2c2f: oData <= 16'h0000;
            14'h2c30: oData <= 16'h0000;
            14'h2c31: oData <= 16'h0000;
            14'h2c32: oData <= 16'h0000;
            14'h2c33: oData <= 16'h0000;
            14'h2c34: oData <= 16'h0000;
            14'h2c35: oData <= 16'h0000;
            14'h2c36: oData <= 16'h0000;
            14'h2c37: oData <= 16'h0000;
            14'h2c38: oData <= 16'h0000;
            14'h2c39: oData <= 16'h0000;
            14'h2c3a: oData <= 16'h0000;
            14'h2c3b: oData <= 16'h0000;
            14'h2c3c: oData <= 16'h0000;
            14'h2c3d: oData <= 16'h0000;
            14'h2c3e: oData <= 16'h0000;
            14'h2c3f: oData <= 16'h0000;
            14'h2c40: oData <= 16'h0000;
            14'h2c41: oData <= 16'h0000;
            14'h2c42: oData <= 16'h0000;
            14'h2c43: oData <= 16'h0000;
            14'h2c44: oData <= 16'h0000;
            14'h2c45: oData <= 16'h0000;
            14'h2c46: oData <= 16'h0000;
            14'h2c47: oData <= 16'h0000;
            14'h2c48: oData <= 16'h0000;
            14'h2c49: oData <= 16'h0000;
            14'h2c4a: oData <= 16'h0000;
            14'h2c4b: oData <= 16'h0000;
            14'h2c4c: oData <= 16'h0000;
            14'h2c4d: oData <= 16'h0000;
            14'h2c4e: oData <= 16'h0000;
            14'h2c4f: oData <= 16'h0000;
            14'h2c50: oData <= 16'h0000;
            14'h2c51: oData <= 16'h0000;
            14'h2c52: oData <= 16'h0000;
            14'h2c53: oData <= 16'h0000;
            14'h2c54: oData <= 16'h0000;
            14'h2c55: oData <= 16'h0000;
            14'h2c56: oData <= 16'h0000;
            14'h2c57: oData <= 16'h0000;
            14'h2c58: oData <= 16'h0000;
            14'h2c59: oData <= 16'h0000;
            14'h2c5a: oData <= 16'h0000;
            14'h2c5b: oData <= 16'h0000;
            14'h2c5c: oData <= 16'h0000;
            14'h2c5d: oData <= 16'h0000;
            14'h2c5e: oData <= 16'h0000;
            14'h2c5f: oData <= 16'h0000;
            14'h2c60: oData <= 16'h0000;
            14'h2c61: oData <= 16'h0000;
            14'h2c62: oData <= 16'h0000;
            14'h2c63: oData <= 16'h0000;
            14'h2c64: oData <= 16'h0000;
            14'h2c65: oData <= 16'h0000;
            14'h2c66: oData <= 16'h0000;
            14'h2c67: oData <= 16'h0000;
            14'h2c68: oData <= 16'h0000;
            14'h2c69: oData <= 16'h0000;
            14'h2c6a: oData <= 16'h0000;
            14'h2c6b: oData <= 16'h0000;
            14'h2c6c: oData <= 16'h0000;
            14'h2c6d: oData <= 16'h0000;
            14'h2c6e: oData <= 16'h0000;
            14'h2c6f: oData <= 16'h0000;
            14'h2c70: oData <= 16'h0000;
            14'h2c71: oData <= 16'h0000;
            14'h2c72: oData <= 16'h0000;
            14'h2c73: oData <= 16'h0000;
            14'h2c74: oData <= 16'h0000;
            14'h2c75: oData <= 16'h0000;
            14'h2c76: oData <= 16'h0000;
            14'h2c77: oData <= 16'h0000;
            14'h2c78: oData <= 16'h0000;
            14'h2c79: oData <= 16'h0000;
            14'h2c7a: oData <= 16'h0000;
            14'h2c7b: oData <= 16'h0000;
            14'h2c7c: oData <= 16'h0000;
            14'h2c7d: oData <= 16'h0000;
            14'h2c7e: oData <= 16'h0000;
            14'h2c7f: oData <= 16'h0000;
            14'h2c80: oData <= 16'h0000;
            14'h2c81: oData <= 16'h0000;
            14'h2c82: oData <= 16'h0000;
            14'h2c83: oData <= 16'h0000;
            14'h2c84: oData <= 16'h0000;
            14'h2c85: oData <= 16'h0000;
            14'h2c86: oData <= 16'h0000;
            14'h2c87: oData <= 16'h0000;
            14'h2c88: oData <= 16'h0000;
            14'h2c89: oData <= 16'h0000;
            14'h2c8a: oData <= 16'h0000;
            14'h2c8b: oData <= 16'h0000;
            14'h2c8c: oData <= 16'h0000;
            14'h2c8d: oData <= 16'h0000;
            14'h2c8e: oData <= 16'h0000;
            14'h2c8f: oData <= 16'h0000;
            14'h2c90: oData <= 16'h0000;
            14'h2c91: oData <= 16'h0000;
            14'h2c92: oData <= 16'h0000;
            14'h2c93: oData <= 16'h0000;
            14'h2c94: oData <= 16'h0000;
            14'h2c95: oData <= 16'h0000;
            14'h2c96: oData <= 16'h0000;
            14'h2c97: oData <= 16'h0000;
            14'h2c98: oData <= 16'h0000;
            14'h2c99: oData <= 16'h0000;
            14'h2c9a: oData <= 16'h0000;
            14'h2c9b: oData <= 16'h0000;
            14'h2c9c: oData <= 16'h0000;
            14'h2c9d: oData <= 16'h0000;
            14'h2c9e: oData <= 16'h0000;
            14'h2c9f: oData <= 16'h0000;
            14'h2ca0: oData <= 16'h0000;
            14'h2ca1: oData <= 16'h0000;
            14'h2ca2: oData <= 16'h0000;
            14'h2ca3: oData <= 16'h0000;
            14'h2ca4: oData <= 16'h0000;
            14'h2ca5: oData <= 16'h0000;
            14'h2ca6: oData <= 16'h0000;
            14'h2ca7: oData <= 16'h0000;
            14'h2ca8: oData <= 16'h0000;
            14'h2ca9: oData <= 16'h0000;
            14'h2caa: oData <= 16'h0000;
            14'h2cab: oData <= 16'h0000;
            14'h2cac: oData <= 16'h0000;
            14'h2cad: oData <= 16'h0000;
            14'h2cae: oData <= 16'h0000;
            14'h2caf: oData <= 16'h0000;
            14'h2cb0: oData <= 16'h0000;
            14'h2cb1: oData <= 16'h0000;
            14'h2cb2: oData <= 16'h0000;
            14'h2cb3: oData <= 16'h0000;
            14'h2cb4: oData <= 16'h0000;
            14'h2cb5: oData <= 16'h0000;
            14'h2cb6: oData <= 16'h0000;
            14'h2cb7: oData <= 16'h0000;
            14'h2cb8: oData <= 16'h0000;
            14'h2cb9: oData <= 16'h0000;
            14'h2cba: oData <= 16'h0000;
            14'h2cbb: oData <= 16'h0000;
            14'h2cbc: oData <= 16'h0000;
            14'h2cbd: oData <= 16'h0000;
            14'h2cbe: oData <= 16'h0000;
            14'h2cbf: oData <= 16'h0000;
            14'h2cc0: oData <= 16'h0000;
            14'h2cc1: oData <= 16'h0000;
            14'h2cc2: oData <= 16'h0000;
            14'h2cc3: oData <= 16'h0000;
            14'h2cc4: oData <= 16'h0000;
            14'h2cc5: oData <= 16'h0000;
            14'h2cc6: oData <= 16'h0000;
            14'h2cc7: oData <= 16'h0000;
            14'h2cc8: oData <= 16'h0000;
            14'h2cc9: oData <= 16'h0000;
            14'h2cca: oData <= 16'h0000;
            14'h2ccb: oData <= 16'h0000;
            14'h2ccc: oData <= 16'h0000;
            14'h2ccd: oData <= 16'h0000;
            14'h2cce: oData <= 16'h0000;
            14'h2ccf: oData <= 16'h0000;
            14'h2cd0: oData <= 16'h0000;
            14'h2cd1: oData <= 16'h0000;
            14'h2cd2: oData <= 16'h0000;
            14'h2cd3: oData <= 16'h0000;
            14'h2cd4: oData <= 16'h0000;
            14'h2cd5: oData <= 16'h0000;
            14'h2cd6: oData <= 16'h0000;
            14'h2cd7: oData <= 16'h0000;
            14'h2cd8: oData <= 16'h0000;
            14'h2cd9: oData <= 16'h0000;
            14'h2cda: oData <= 16'h0000;
            14'h2cdb: oData <= 16'h0000;
            14'h2cdc: oData <= 16'h0000;
            14'h2cdd: oData <= 16'h0000;
            14'h2cde: oData <= 16'h0000;
            14'h2cdf: oData <= 16'h0000;
            14'h2ce0: oData <= 16'h0000;
            14'h2ce1: oData <= 16'h0000;
            14'h2ce2: oData <= 16'h0000;
            14'h2ce3: oData <= 16'h0000;
            14'h2ce4: oData <= 16'h0000;
            14'h2ce5: oData <= 16'h0000;
            14'h2ce6: oData <= 16'h0000;
            14'h2ce7: oData <= 16'h0000;
            14'h2ce8: oData <= 16'h0000;
            14'h2ce9: oData <= 16'h0000;
            14'h2cea: oData <= 16'h0000;
            14'h2ceb: oData <= 16'h0000;
            14'h2cec: oData <= 16'h0000;
            14'h2ced: oData <= 16'h0000;
            14'h2cee: oData <= 16'h0000;
            14'h2cef: oData <= 16'h0000;
            14'h2cf0: oData <= 16'h0000;
            14'h2cf1: oData <= 16'h0000;
            14'h2cf2: oData <= 16'h0000;
            14'h2cf3: oData <= 16'h0000;
            14'h2cf4: oData <= 16'h0000;
            14'h2cf5: oData <= 16'h0000;
            14'h2cf6: oData <= 16'h0000;
            14'h2cf7: oData <= 16'h0000;
            14'h2cf8: oData <= 16'h0000;
            14'h2cf9: oData <= 16'h0000;
            14'h2cfa: oData <= 16'h0000;
            14'h2cfb: oData <= 16'h0000;
            14'h2cfc: oData <= 16'h0000;
            14'h2cfd: oData <= 16'h0000;
            14'h2cfe: oData <= 16'h0000;
            14'h2cff: oData <= 16'h0000;
            14'h2d00: oData <= 16'h0000;
            14'h2d01: oData <= 16'h0000;
            14'h2d02: oData <= 16'h0000;
            14'h2d03: oData <= 16'h0000;
            14'h2d04: oData <= 16'h0000;
            14'h2d05: oData <= 16'h0000;
            14'h2d06: oData <= 16'h0000;
            14'h2d07: oData <= 16'h0000;
            14'h2d08: oData <= 16'h0000;
            14'h2d09: oData <= 16'h0000;
            14'h2d0a: oData <= 16'h0000;
            14'h2d0b: oData <= 16'h0000;
            14'h2d0c: oData <= 16'h0000;
            14'h2d0d: oData <= 16'h0000;
            14'h2d0e: oData <= 16'h0000;
            14'h2d0f: oData <= 16'h0000;
            14'h2d10: oData <= 16'h0000;
            14'h2d11: oData <= 16'h0000;
            14'h2d12: oData <= 16'h0000;
            14'h2d13: oData <= 16'h0000;
            14'h2d14: oData <= 16'h0000;
            14'h2d15: oData <= 16'h0000;
            14'h2d16: oData <= 16'h0000;
            14'h2d17: oData <= 16'h0000;
            14'h2d18: oData <= 16'h0000;
            14'h2d19: oData <= 16'h0000;
            14'h2d1a: oData <= 16'h0000;
            14'h2d1b: oData <= 16'h0000;
            14'h2d1c: oData <= 16'h0000;
            14'h2d1d: oData <= 16'h0000;
            14'h2d1e: oData <= 16'h0000;
            14'h2d1f: oData <= 16'h0000;
            14'h2d20: oData <= 16'h0000;
            14'h2d21: oData <= 16'h0000;
            14'h2d22: oData <= 16'h0000;
            14'h2d23: oData <= 16'h0000;
            14'h2d24: oData <= 16'h0000;
            14'h2d25: oData <= 16'h0000;
            14'h2d26: oData <= 16'h0000;
            14'h2d27: oData <= 16'h0000;
            14'h2d28: oData <= 16'h0000;
            14'h2d29: oData <= 16'h0000;
            14'h2d2a: oData <= 16'h0000;
            14'h2d2b: oData <= 16'h0000;
            14'h2d2c: oData <= 16'h0000;
            14'h2d2d: oData <= 16'h0000;
            14'h2d2e: oData <= 16'h0000;
            14'h2d2f: oData <= 16'h0000;
            14'h2d30: oData <= 16'h0000;
            14'h2d31: oData <= 16'h0000;
            14'h2d32: oData <= 16'h0000;
            14'h2d33: oData <= 16'h0000;
            14'h2d34: oData <= 16'h0000;
            14'h2d35: oData <= 16'h0000;
            14'h2d36: oData <= 16'h0000;
            14'h2d37: oData <= 16'h0000;
            14'h2d38: oData <= 16'h0000;
            14'h2d39: oData <= 16'h0000;
            14'h2d3a: oData <= 16'h0000;
            14'h2d3b: oData <= 16'h0000;
            14'h2d3c: oData <= 16'h0000;
            14'h2d3d: oData <= 16'h0000;
            14'h2d3e: oData <= 16'h0000;
            14'h2d3f: oData <= 16'h0000;
            14'h2d40: oData <= 16'h0000;
            14'h2d41: oData <= 16'h0000;
            14'h2d42: oData <= 16'h0000;
            14'h2d43: oData <= 16'h0000;
            14'h2d44: oData <= 16'h0000;
            14'h2d45: oData <= 16'h0000;
            14'h2d46: oData <= 16'h0000;
            14'h2d47: oData <= 16'h0000;
            14'h2d48: oData <= 16'h0000;
            14'h2d49: oData <= 16'h0000;
            14'h2d4a: oData <= 16'h0000;
            14'h2d4b: oData <= 16'h0000;
            14'h2d4c: oData <= 16'h0000;
            14'h2d4d: oData <= 16'h0000;
            14'h2d4e: oData <= 16'h0000;
            14'h2d4f: oData <= 16'h0000;
            14'h2d50: oData <= 16'h0000;
            14'h2d51: oData <= 16'h0000;
            14'h2d52: oData <= 16'h0000;
            14'h2d53: oData <= 16'h0000;
            14'h2d54: oData <= 16'h0000;
            14'h2d55: oData <= 16'h0000;
            14'h2d56: oData <= 16'h0000;
            14'h2d57: oData <= 16'h0000;
            14'h2d58: oData <= 16'h0000;
            14'h2d59: oData <= 16'h0000;
            14'h2d5a: oData <= 16'h0000;
            14'h2d5b: oData <= 16'h0000;
            14'h2d5c: oData <= 16'h0000;
            14'h2d5d: oData <= 16'h0000;
            14'h2d5e: oData <= 16'h0000;
            14'h2d5f: oData <= 16'h0000;
            14'h2d60: oData <= 16'h0000;
            14'h2d61: oData <= 16'h0000;
            14'h2d62: oData <= 16'h0000;
            14'h2d63: oData <= 16'h0000;
            14'h2d64: oData <= 16'h0000;
            14'h2d65: oData <= 16'h0000;
            14'h2d66: oData <= 16'h0000;
            14'h2d67: oData <= 16'h0000;
            14'h2d68: oData <= 16'h0000;
            14'h2d69: oData <= 16'h0000;
            14'h2d6a: oData <= 16'h0000;
            14'h2d6b: oData <= 16'h0000;
            14'h2d6c: oData <= 16'h0000;
            14'h2d6d: oData <= 16'h0000;
            14'h2d6e: oData <= 16'h0000;
            14'h2d6f: oData <= 16'h0000;
            14'h2d70: oData <= 16'h0000;
            14'h2d71: oData <= 16'h0000;
            14'h2d72: oData <= 16'h0000;
            14'h2d73: oData <= 16'h0000;
            14'h2d74: oData <= 16'h0000;
            14'h2d75: oData <= 16'h0000;
            14'h2d76: oData <= 16'h0000;
            14'h2d77: oData <= 16'h0000;
            14'h2d78: oData <= 16'h0000;
            14'h2d79: oData <= 16'h0000;
            14'h2d7a: oData <= 16'h0000;
            14'h2d7b: oData <= 16'h0000;
            14'h2d7c: oData <= 16'h0000;
            14'h2d7d: oData <= 16'h0000;
            14'h2d7e: oData <= 16'h0000;
            14'h2d7f: oData <= 16'h0000;
            14'h2d80: oData <= 16'h0000;
            14'h2d81: oData <= 16'h0000;
            14'h2d82: oData <= 16'h0000;
            14'h2d83: oData <= 16'h0000;
            14'h2d84: oData <= 16'h0000;
            14'h2d85: oData <= 16'h0000;
            14'h2d86: oData <= 16'h0000;
            14'h2d87: oData <= 16'h0000;
            14'h2d88: oData <= 16'h0000;
            14'h2d89: oData <= 16'h0000;
            14'h2d8a: oData <= 16'h0000;
            14'h2d8b: oData <= 16'h0000;
            14'h2d8c: oData <= 16'h0000;
            14'h2d8d: oData <= 16'h0000;
            14'h2d8e: oData <= 16'h0000;
            14'h2d8f: oData <= 16'h0000;
            14'h2d90: oData <= 16'h0000;
            14'h2d91: oData <= 16'h0000;
            14'h2d92: oData <= 16'h0000;
            14'h2d93: oData <= 16'h0000;
            14'h2d94: oData <= 16'h0000;
            14'h2d95: oData <= 16'h0000;
            14'h2d96: oData <= 16'h0000;
            14'h2d97: oData <= 16'h0000;
            14'h2d98: oData <= 16'h0000;
            14'h2d99: oData <= 16'h0000;
            14'h2d9a: oData <= 16'h0000;
            14'h2d9b: oData <= 16'h0000;
            14'h2d9c: oData <= 16'h0000;
            14'h2d9d: oData <= 16'h0000;
            14'h2d9e: oData <= 16'h0000;
            14'h2d9f: oData <= 16'h0000;
            14'h2da0: oData <= 16'h0000;
            14'h2da1: oData <= 16'h0000;
            14'h2da2: oData <= 16'h0000;
            14'h2da3: oData <= 16'h0000;
            14'h2da4: oData <= 16'h0000;
            14'h2da5: oData <= 16'h0000;
            14'h2da6: oData <= 16'h0000;
            14'h2da7: oData <= 16'h0000;
            14'h2da8: oData <= 16'h0000;
            14'h2da9: oData <= 16'h0000;
            14'h2daa: oData <= 16'h0000;
            14'h2dab: oData <= 16'h0000;
            14'h2dac: oData <= 16'h0000;
            14'h2dad: oData <= 16'h0000;
            14'h2dae: oData <= 16'h0000;
            14'h2daf: oData <= 16'h0000;
            14'h2db0: oData <= 16'h0000;
            14'h2db1: oData <= 16'h0000;
            14'h2db2: oData <= 16'h0000;
            14'h2db3: oData <= 16'h0000;
            14'h2db4: oData <= 16'h0000;
            14'h2db5: oData <= 16'h0000;
            14'h2db6: oData <= 16'h0000;
            14'h2db7: oData <= 16'h0000;
            14'h2db8: oData <= 16'h0000;
            14'h2db9: oData <= 16'h0000;
            14'h2dba: oData <= 16'h0000;
            14'h2dbb: oData <= 16'h0000;
            14'h2dbc: oData <= 16'h0000;
            14'h2dbd: oData <= 16'h0000;
            14'h2dbe: oData <= 16'h0000;
            14'h2dbf: oData <= 16'h0000;
            14'h2dc0: oData <= 16'h0000;
            14'h2dc1: oData <= 16'h0000;
            14'h2dc2: oData <= 16'h0000;
            14'h2dc3: oData <= 16'h0000;
            14'h2dc4: oData <= 16'h0000;
            14'h2dc5: oData <= 16'h0000;
            14'h2dc6: oData <= 16'h0000;
            14'h2dc7: oData <= 16'h0000;
            14'h2dc8: oData <= 16'h0000;
            14'h2dc9: oData <= 16'h0000;
            14'h2dca: oData <= 16'h0000;
            14'h2dcb: oData <= 16'h0000;
            14'h2dcc: oData <= 16'h0000;
            14'h2dcd: oData <= 16'h0000;
            14'h2dce: oData <= 16'h0000;
            14'h2dcf: oData <= 16'h0000;
            14'h2dd0: oData <= 16'h0000;
            14'h2dd1: oData <= 16'h0000;
            14'h2dd2: oData <= 16'h0000;
            14'h2dd3: oData <= 16'h0000;
            14'h2dd4: oData <= 16'h0000;
            14'h2dd5: oData <= 16'h0000;
            14'h2dd6: oData <= 16'h0000;
            14'h2dd7: oData <= 16'h0000;
            14'h2dd8: oData <= 16'h0000;
            14'h2dd9: oData <= 16'h0000;
            14'h2dda: oData <= 16'h0000;
            14'h2ddb: oData <= 16'h0000;
            14'h2ddc: oData <= 16'h0000;
            14'h2ddd: oData <= 16'h0000;
            14'h2dde: oData <= 16'h0000;
            14'h2ddf: oData <= 16'h0000;
            14'h2de0: oData <= 16'h0000;
            14'h2de1: oData <= 16'h0000;
            14'h2de2: oData <= 16'h0000;
            14'h2de3: oData <= 16'h0000;
            14'h2de4: oData <= 16'h0000;
            14'h2de5: oData <= 16'h0000;
            14'h2de6: oData <= 16'h0000;
            14'h2de7: oData <= 16'h0000;
            14'h2de8: oData <= 16'h0000;
            14'h2de9: oData <= 16'h0000;
            14'h2dea: oData <= 16'h0000;
            14'h2deb: oData <= 16'h0000;
            14'h2dec: oData <= 16'h0000;
            14'h2ded: oData <= 16'h0000;
            14'h2dee: oData <= 16'h0000;
            14'h2def: oData <= 16'h0000;
            14'h2df0: oData <= 16'h0000;
            14'h2df1: oData <= 16'h0000;
            14'h2df2: oData <= 16'h0000;
            14'h2df3: oData <= 16'h0000;
            14'h2df4: oData <= 16'h0000;
            14'h2df5: oData <= 16'h0000;
            14'h2df6: oData <= 16'h0000;
            14'h2df7: oData <= 16'h0000;
            14'h2df8: oData <= 16'h0000;
            14'h2df9: oData <= 16'h0000;
            14'h2dfa: oData <= 16'h0000;
            14'h2dfb: oData <= 16'h0000;
            14'h2dfc: oData <= 16'h0000;
            14'h2dfd: oData <= 16'h0000;
            14'h2dfe: oData <= 16'h0000;
            14'h2dff: oData <= 16'h0000;
            14'h2e00: oData <= 16'h0000;
            14'h2e01: oData <= 16'h0000;
            14'h2e02: oData <= 16'h0000;
            14'h2e03: oData <= 16'h0000;
            14'h2e04: oData <= 16'h0000;
            14'h2e05: oData <= 16'h0000;
            14'h2e06: oData <= 16'h0000;
            14'h2e07: oData <= 16'h0000;
            14'h2e08: oData <= 16'h0000;
            14'h2e09: oData <= 16'h0000;
            14'h2e0a: oData <= 16'h0000;
            14'h2e0b: oData <= 16'h0000;
            14'h2e0c: oData <= 16'h0000;
            14'h2e0d: oData <= 16'h0000;
            14'h2e0e: oData <= 16'h0000;
            14'h2e0f: oData <= 16'h0000;
            14'h2e10: oData <= 16'h0000;
            14'h2e11: oData <= 16'h0000;
            14'h2e12: oData <= 16'h0000;
            14'h2e13: oData <= 16'h0000;
            14'h2e14: oData <= 16'h0000;
            14'h2e15: oData <= 16'h0000;
            14'h2e16: oData <= 16'h0000;
            14'h2e17: oData <= 16'h0000;
            14'h2e18: oData <= 16'h0000;
            14'h2e19: oData <= 16'h0000;
            14'h2e1a: oData <= 16'h0000;
            14'h2e1b: oData <= 16'h0000;
            14'h2e1c: oData <= 16'h0000;
            14'h2e1d: oData <= 16'h0000;
            14'h2e1e: oData <= 16'h0000;
            14'h2e1f: oData <= 16'h0000;
            14'h2e20: oData <= 16'h0000;
            14'h2e21: oData <= 16'h0000;
            14'h2e22: oData <= 16'h0000;
            14'h2e23: oData <= 16'h0000;
            14'h2e24: oData <= 16'h0000;
            14'h2e25: oData <= 16'h0000;
            14'h2e26: oData <= 16'h0000;
            14'h2e27: oData <= 16'h0000;
            14'h2e28: oData <= 16'h0000;
            14'h2e29: oData <= 16'h0000;
            14'h2e2a: oData <= 16'h0000;
            14'h2e2b: oData <= 16'h0000;
            14'h2e2c: oData <= 16'h0000;
            14'h2e2d: oData <= 16'h0000;
            14'h2e2e: oData <= 16'h0000;
            14'h2e2f: oData <= 16'h0000;
            14'h2e30: oData <= 16'h0000;
            14'h2e31: oData <= 16'h0000;
            14'h2e32: oData <= 16'h0000;
            14'h2e33: oData <= 16'h0000;
            14'h2e34: oData <= 16'h0000;
            14'h2e35: oData <= 16'h0000;
            14'h2e36: oData <= 16'h0000;
            14'h2e37: oData <= 16'h0000;
            14'h2e38: oData <= 16'h0000;
            14'h2e39: oData <= 16'h0000;
            14'h2e3a: oData <= 16'h0000;
            14'h2e3b: oData <= 16'h0000;
            14'h2e3c: oData <= 16'h0000;
            14'h2e3d: oData <= 16'h0000;
            14'h2e3e: oData <= 16'h0000;
            14'h2e3f: oData <= 16'h0000;
            14'h2e40: oData <= 16'h0000;
            14'h2e41: oData <= 16'h0000;
            14'h2e42: oData <= 16'h0000;
            14'h2e43: oData <= 16'h0000;
            14'h2e44: oData <= 16'h0000;
            14'h2e45: oData <= 16'h0000;
            14'h2e46: oData <= 16'h0000;
            14'h2e47: oData <= 16'h0000;
            14'h2e48: oData <= 16'h0000;
            14'h2e49: oData <= 16'h0000;
            14'h2e4a: oData <= 16'h0000;
            14'h2e4b: oData <= 16'h0000;
            14'h2e4c: oData <= 16'h0000;
            14'h2e4d: oData <= 16'h0000;
            14'h2e4e: oData <= 16'h0000;
            14'h2e4f: oData <= 16'h0000;
            14'h2e50: oData <= 16'h0000;
            14'h2e51: oData <= 16'h0000;
            14'h2e52: oData <= 16'h0000;
            14'h2e53: oData <= 16'h0000;
            14'h2e54: oData <= 16'h0000;
            14'h2e55: oData <= 16'h0000;
            14'h2e56: oData <= 16'h0000;
            14'h2e57: oData <= 16'h0000;
            14'h2e58: oData <= 16'h0000;
            14'h2e59: oData <= 16'h0000;
            14'h2e5a: oData <= 16'h0000;
            14'h2e5b: oData <= 16'h0000;
            14'h2e5c: oData <= 16'h0000;
            14'h2e5d: oData <= 16'h0000;
            14'h2e5e: oData <= 16'h0000;
            14'h2e5f: oData <= 16'h0000;
            14'h2e60: oData <= 16'h0000;
            14'h2e61: oData <= 16'h0000;
            14'h2e62: oData <= 16'h0000;
            14'h2e63: oData <= 16'h0000;
            14'h2e64: oData <= 16'h0000;
            14'h2e65: oData <= 16'h0000;
            14'h2e66: oData <= 16'h0000;
            14'h2e67: oData <= 16'h0000;
            14'h2e68: oData <= 16'h0000;
            14'h2e69: oData <= 16'h0000;
            14'h2e6a: oData <= 16'h0000;
            14'h2e6b: oData <= 16'h0000;
            14'h2e6c: oData <= 16'h0000;
            14'h2e6d: oData <= 16'h0000;
            14'h2e6e: oData <= 16'h0000;
            14'h2e6f: oData <= 16'h0000;
            14'h2e70: oData <= 16'h0000;
            14'h2e71: oData <= 16'h0000;
            14'h2e72: oData <= 16'h0000;
            14'h2e73: oData <= 16'h0000;
            14'h2e74: oData <= 16'h0000;
            14'h2e75: oData <= 16'h0000;
            14'h2e76: oData <= 16'h0000;
            14'h2e77: oData <= 16'h0000;
            14'h2e78: oData <= 16'h0000;
            14'h2e79: oData <= 16'h0000;
            14'h2e7a: oData <= 16'h0000;
            14'h2e7b: oData <= 16'h0000;
            14'h2e7c: oData <= 16'h0000;
            14'h2e7d: oData <= 16'h0000;
            14'h2e7e: oData <= 16'h0000;
            14'h2e7f: oData <= 16'h0000;
            14'h2e80: oData <= 16'h0000;
            14'h2e81: oData <= 16'h0000;
            14'h2e82: oData <= 16'h0000;
            14'h2e83: oData <= 16'h0000;
            14'h2e84: oData <= 16'h0000;
            14'h2e85: oData <= 16'h0000;
            14'h2e86: oData <= 16'h0000;
            14'h2e87: oData <= 16'h0000;
            14'h2e88: oData <= 16'h0000;
            14'h2e89: oData <= 16'h0000;
            14'h2e8a: oData <= 16'h0000;
            14'h2e8b: oData <= 16'h0000;
            14'h2e8c: oData <= 16'h0000;
            14'h2e8d: oData <= 16'h0000;
            14'h2e8e: oData <= 16'h0000;
            14'h2e8f: oData <= 16'h0000;
            14'h2e90: oData <= 16'h0000;
            14'h2e91: oData <= 16'h0000;
            14'h2e92: oData <= 16'h0000;
            14'h2e93: oData <= 16'h0000;
            14'h2e94: oData <= 16'h0000;
            14'h2e95: oData <= 16'h0000;
            14'h2e96: oData <= 16'h0000;
            14'h2e97: oData <= 16'h0000;
            14'h2e98: oData <= 16'h0000;
            14'h2e99: oData <= 16'h0000;
            14'h2e9a: oData <= 16'h0000;
            14'h2e9b: oData <= 16'h0000;
            14'h2e9c: oData <= 16'h0000;
            14'h2e9d: oData <= 16'h0000;
            14'h2e9e: oData <= 16'h0000;
            14'h2e9f: oData <= 16'h0000;
            14'h2ea0: oData <= 16'h0000;
            14'h2ea1: oData <= 16'h0000;
            14'h2ea2: oData <= 16'h0000;
            14'h2ea3: oData <= 16'h0000;
            14'h2ea4: oData <= 16'h0000;
            14'h2ea5: oData <= 16'h0000;
            14'h2ea6: oData <= 16'h0000;
            14'h2ea7: oData <= 16'h0000;
            14'h2ea8: oData <= 16'h0000;
            14'h2ea9: oData <= 16'h0000;
            14'h2eaa: oData <= 16'h0000;
            14'h2eab: oData <= 16'h0000;
            14'h2eac: oData <= 16'h0000;
            14'h2ead: oData <= 16'h0000;
            14'h2eae: oData <= 16'h0000;
            14'h2eaf: oData <= 16'h0000;
            14'h2eb0: oData <= 16'h0000;
            14'h2eb1: oData <= 16'h0000;
            14'h2eb2: oData <= 16'h0000;
            14'h2eb3: oData <= 16'h0000;
            14'h2eb4: oData <= 16'h0000;
            14'h2eb5: oData <= 16'h0000;
            14'h2eb6: oData <= 16'h0000;
            14'h2eb7: oData <= 16'h0000;
            14'h2eb8: oData <= 16'h0000;
            14'h2eb9: oData <= 16'h0000;
            14'h2eba: oData <= 16'h0000;
            14'h2ebb: oData <= 16'h0000;
            14'h2ebc: oData <= 16'h0000;
            14'h2ebd: oData <= 16'h0000;
            14'h2ebe: oData <= 16'h0000;
            14'h2ebf: oData <= 16'h0000;
            14'h2ec0: oData <= 16'h0000;
            14'h2ec1: oData <= 16'h0000;
            14'h2ec2: oData <= 16'h0000;
            14'h2ec3: oData <= 16'h0000;
            14'h2ec4: oData <= 16'h0000;
            14'h2ec5: oData <= 16'h0000;
            14'h2ec6: oData <= 16'h0000;
            14'h2ec7: oData <= 16'h0000;
            14'h2ec8: oData <= 16'h0000;
            14'h2ec9: oData <= 16'h0000;
            14'h2eca: oData <= 16'h0000;
            14'h2ecb: oData <= 16'h0000;
            14'h2ecc: oData <= 16'h0000;
            14'h2ecd: oData <= 16'h0000;
            14'h2ece: oData <= 16'h0000;
            14'h2ecf: oData <= 16'h0000;
            14'h2ed0: oData <= 16'h0000;
            14'h2ed1: oData <= 16'h0000;
            14'h2ed2: oData <= 16'h0000;
            14'h2ed3: oData <= 16'h0000;
            14'h2ed4: oData <= 16'h0000;
            14'h2ed5: oData <= 16'h0000;
            14'h2ed6: oData <= 16'h0000;
            14'h2ed7: oData <= 16'h0000;
            14'h2ed8: oData <= 16'h0000;
            14'h2ed9: oData <= 16'h0000;
            14'h2eda: oData <= 16'h0000;
            14'h2edb: oData <= 16'h0000;
            14'h2edc: oData <= 16'h0000;
            14'h2edd: oData <= 16'h0000;
            14'h2ede: oData <= 16'h0000;
            14'h2edf: oData <= 16'h0000;
            14'h2ee0: oData <= 16'h0000;
            14'h2ee1: oData <= 16'h0000;
            14'h2ee2: oData <= 16'h0000;
            14'h2ee3: oData <= 16'h0000;
            14'h2ee4: oData <= 16'h0000;
            14'h2ee5: oData <= 16'h0000;
            14'h2ee6: oData <= 16'h0000;
            14'h2ee7: oData <= 16'h0000;
            14'h2ee8: oData <= 16'h0000;
            14'h2ee9: oData <= 16'h0000;
            14'h2eea: oData <= 16'h0000;
            14'h2eeb: oData <= 16'h0000;
            14'h2eec: oData <= 16'h0000;
            14'h2eed: oData <= 16'h0000;
            14'h2eee: oData <= 16'h0000;
            14'h2eef: oData <= 16'h0000;
            14'h2ef0: oData <= 16'h0000;
            14'h2ef1: oData <= 16'h0000;
            14'h2ef2: oData <= 16'h0000;
            14'h2ef3: oData <= 16'h0000;
            14'h2ef4: oData <= 16'h0000;
            14'h2ef5: oData <= 16'h0000;
            14'h2ef6: oData <= 16'h0000;
            14'h2ef7: oData <= 16'h0000;
            14'h2ef8: oData <= 16'h0000;
            14'h2ef9: oData <= 16'h0000;
            14'h2efa: oData <= 16'h0000;
            14'h2efb: oData <= 16'h0000;
            14'h2efc: oData <= 16'h0000;
            14'h2efd: oData <= 16'h0000;
            14'h2efe: oData <= 16'h0000;
            14'h2eff: oData <= 16'h0000;
            14'h2f00: oData <= 16'h0000;
            14'h2f01: oData <= 16'h0000;
            14'h2f02: oData <= 16'h0000;
            14'h2f03: oData <= 16'h0000;
            14'h2f04: oData <= 16'h0000;
            14'h2f05: oData <= 16'h0000;
            14'h2f06: oData <= 16'h0000;
            14'h2f07: oData <= 16'h0000;
            14'h2f08: oData <= 16'h0000;
            14'h2f09: oData <= 16'h0000;
            14'h2f0a: oData <= 16'h0000;
            14'h2f0b: oData <= 16'h0000;
            14'h2f0c: oData <= 16'h0000;
            14'h2f0d: oData <= 16'h0000;
            14'h2f0e: oData <= 16'h0000;
            14'h2f0f: oData <= 16'h0000;
            14'h2f10: oData <= 16'h0000;
            14'h2f11: oData <= 16'h0000;
            14'h2f12: oData <= 16'h0000;
            14'h2f13: oData <= 16'h0000;
            14'h2f14: oData <= 16'h0000;
            14'h2f15: oData <= 16'h0000;
            14'h2f16: oData <= 16'h0000;
            14'h2f17: oData <= 16'h0000;
            14'h2f18: oData <= 16'h0000;
            14'h2f19: oData <= 16'h0000;
            14'h2f1a: oData <= 16'h0000;
            14'h2f1b: oData <= 16'h0000;
            14'h2f1c: oData <= 16'h0000;
            14'h2f1d: oData <= 16'h0000;
            14'h2f1e: oData <= 16'h0000;
            14'h2f1f: oData <= 16'h0000;
            14'h2f20: oData <= 16'h0000;
            14'h2f21: oData <= 16'h0000;
            14'h2f22: oData <= 16'h0000;
            14'h2f23: oData <= 16'h0000;
            14'h2f24: oData <= 16'h0000;
            14'h2f25: oData <= 16'h0000;
            14'h2f26: oData <= 16'h0000;
            14'h2f27: oData <= 16'h0000;
            14'h2f28: oData <= 16'h0000;
            14'h2f29: oData <= 16'h0000;
            14'h2f2a: oData <= 16'h0000;
            14'h2f2b: oData <= 16'h0000;
            14'h2f2c: oData <= 16'h0000;
            14'h2f2d: oData <= 16'h0000;
            14'h2f2e: oData <= 16'h0000;
            14'h2f2f: oData <= 16'h0000;
            14'h2f30: oData <= 16'h0000;
            14'h2f31: oData <= 16'h0000;
            14'h2f32: oData <= 16'h0000;
            14'h2f33: oData <= 16'h0000;
            14'h2f34: oData <= 16'h0000;
            14'h2f35: oData <= 16'h0000;
            14'h2f36: oData <= 16'h0000;
            14'h2f37: oData <= 16'h0000;
            14'h2f38: oData <= 16'h0000;
            14'h2f39: oData <= 16'h0000;
            14'h2f3a: oData <= 16'h0000;
            14'h2f3b: oData <= 16'h0000;
            14'h2f3c: oData <= 16'h0000;
            14'h2f3d: oData <= 16'h0000;
            14'h2f3e: oData <= 16'h0000;
            14'h2f3f: oData <= 16'h0000;
            14'h2f40: oData <= 16'h0000;
            14'h2f41: oData <= 16'h0000;
            14'h2f42: oData <= 16'h0000;
            14'h2f43: oData <= 16'h0000;
            14'h2f44: oData <= 16'h0000;
            14'h2f45: oData <= 16'h0000;
            14'h2f46: oData <= 16'h0000;
            14'h2f47: oData <= 16'h0000;
            14'h2f48: oData <= 16'h0000;
            14'h2f49: oData <= 16'h0000;
            14'h2f4a: oData <= 16'h0000;
            14'h2f4b: oData <= 16'h0000;
            14'h2f4c: oData <= 16'h0000;
            14'h2f4d: oData <= 16'h0000;
            14'h2f4e: oData <= 16'h0000;
            14'h2f4f: oData <= 16'h0000;
            14'h2f50: oData <= 16'h0000;
            14'h2f51: oData <= 16'h0000;
            14'h2f52: oData <= 16'h0000;
            14'h2f53: oData <= 16'h0000;
            14'h2f54: oData <= 16'h0000;
            14'h2f55: oData <= 16'h0000;
            14'h2f56: oData <= 16'h0000;
            14'h2f57: oData <= 16'h0000;
            14'h2f58: oData <= 16'h0000;
            14'h2f59: oData <= 16'h0000;
            14'h2f5a: oData <= 16'h0000;
            14'h2f5b: oData <= 16'h0000;
            14'h2f5c: oData <= 16'h0000;
            14'h2f5d: oData <= 16'h0000;
            14'h2f5e: oData <= 16'h0000;
            14'h2f5f: oData <= 16'h0000;
            14'h2f60: oData <= 16'h0000;
            14'h2f61: oData <= 16'h0000;
            14'h2f62: oData <= 16'h0000;
            14'h2f63: oData <= 16'h0000;
            14'h2f64: oData <= 16'h0000;
            14'h2f65: oData <= 16'h0000;
            14'h2f66: oData <= 16'h0000;
            14'h2f67: oData <= 16'h0000;
            14'h2f68: oData <= 16'h0000;
            14'h2f69: oData <= 16'h0000;
            14'h2f6a: oData <= 16'h0000;
            14'h2f6b: oData <= 16'h0000;
            14'h2f6c: oData <= 16'h0000;
            14'h2f6d: oData <= 16'h0000;
            14'h2f6e: oData <= 16'h0000;
            14'h2f6f: oData <= 16'h0000;
            14'h2f70: oData <= 16'h0000;
            14'h2f71: oData <= 16'h0000;
            14'h2f72: oData <= 16'h0000;
            14'h2f73: oData <= 16'h0000;
            14'h2f74: oData <= 16'h0000;
            14'h2f75: oData <= 16'h0000;
            14'h2f76: oData <= 16'h0000;
            14'h2f77: oData <= 16'h0000;
            14'h2f78: oData <= 16'h0000;
            14'h2f79: oData <= 16'h0000;
            14'h2f7a: oData <= 16'h0000;
            14'h2f7b: oData <= 16'h0000;
            14'h2f7c: oData <= 16'h0000;
            14'h2f7d: oData <= 16'h0000;
            14'h2f7e: oData <= 16'h0000;
            14'h2f7f: oData <= 16'h0000;
            14'h2f80: oData <= 16'h0000;
            14'h2f81: oData <= 16'h0000;
            14'h2f82: oData <= 16'h0000;
            14'h2f83: oData <= 16'h0000;
            14'h2f84: oData <= 16'h0000;
            14'h2f85: oData <= 16'h0000;
            14'h2f86: oData <= 16'h0000;
            14'h2f87: oData <= 16'h0000;
            14'h2f88: oData <= 16'h0000;
            14'h2f89: oData <= 16'h0000;
            14'h2f8a: oData <= 16'h0000;
            14'h2f8b: oData <= 16'h0000;
            14'h2f8c: oData <= 16'h0000;
            14'h2f8d: oData <= 16'h0000;
            14'h2f8e: oData <= 16'h0000;
            14'h2f8f: oData <= 16'h0000;
            14'h2f90: oData <= 16'h0000;
            14'h2f91: oData <= 16'h0000;
            14'h2f92: oData <= 16'h0000;
            14'h2f93: oData <= 16'h0000;
            14'h2f94: oData <= 16'h0000;
            14'h2f95: oData <= 16'h0000;
            14'h2f96: oData <= 16'h0000;
            14'h2f97: oData <= 16'h0000;
            14'h2f98: oData <= 16'h0000;
            14'h2f99: oData <= 16'h0000;
            14'h2f9a: oData <= 16'h0000;
            14'h2f9b: oData <= 16'h0000;
            14'h2f9c: oData <= 16'h0000;
            14'h2f9d: oData <= 16'h0000;
            14'h2f9e: oData <= 16'h0000;
            14'h2f9f: oData <= 16'h0000;
            14'h2fa0: oData <= 16'h0000;
            14'h2fa1: oData <= 16'h0000;
            14'h2fa2: oData <= 16'h0000;
            14'h2fa3: oData <= 16'h0000;
            14'h2fa4: oData <= 16'h0000;
            14'h2fa5: oData <= 16'h0000;
            14'h2fa6: oData <= 16'h0000;
            14'h2fa7: oData <= 16'h0000;
            14'h2fa8: oData <= 16'h0000;
            14'h2fa9: oData <= 16'h0000;
            14'h2faa: oData <= 16'h0000;
            14'h2fab: oData <= 16'h0000;
            14'h2fac: oData <= 16'h0000;
            14'h2fad: oData <= 16'h0000;
            14'h2fae: oData <= 16'h0000;
            14'h2faf: oData <= 16'h0000;
            14'h2fb0: oData <= 16'h0000;
            14'h2fb1: oData <= 16'h0000;
            14'h2fb2: oData <= 16'h0000;
            14'h2fb3: oData <= 16'h0000;
            14'h2fb4: oData <= 16'h0000;
            14'h2fb5: oData <= 16'h0000;
            14'h2fb6: oData <= 16'h0000;
            14'h2fb7: oData <= 16'h0000;
            14'h2fb8: oData <= 16'h0000;
            14'h2fb9: oData <= 16'h0000;
            14'h2fba: oData <= 16'h0000;
            14'h2fbb: oData <= 16'h0000;
            14'h2fbc: oData <= 16'h0000;
            14'h2fbd: oData <= 16'h0000;
            14'h2fbe: oData <= 16'h0000;
            14'h2fbf: oData <= 16'h0000;
            14'h2fc0: oData <= 16'h0000;
            14'h2fc1: oData <= 16'h0000;
            14'h2fc2: oData <= 16'h0000;
            14'h2fc3: oData <= 16'h0000;
            14'h2fc4: oData <= 16'h0000;
            14'h2fc5: oData <= 16'h0000;
            14'h2fc6: oData <= 16'h0000;
            14'h2fc7: oData <= 16'h0000;
            14'h2fc8: oData <= 16'h0000;
            14'h2fc9: oData <= 16'h0000;
            14'h2fca: oData <= 16'h0000;
            14'h2fcb: oData <= 16'h0000;
            14'h2fcc: oData <= 16'h0000;
            14'h2fcd: oData <= 16'h0000;
            14'h2fce: oData <= 16'h0000;
            14'h2fcf: oData <= 16'h0000;
            14'h2fd0: oData <= 16'h0000;
            14'h2fd1: oData <= 16'h0000;
            14'h2fd2: oData <= 16'h0000;
            14'h2fd3: oData <= 16'h0000;
            14'h2fd4: oData <= 16'h0000;
            14'h2fd5: oData <= 16'h0000;
            14'h2fd6: oData <= 16'h0000;
            14'h2fd7: oData <= 16'h0000;
            14'h2fd8: oData <= 16'h0000;
            14'h2fd9: oData <= 16'h0000;
            14'h2fda: oData <= 16'h0000;
            14'h2fdb: oData <= 16'h0000;
            14'h2fdc: oData <= 16'h0000;
            14'h2fdd: oData <= 16'h0000;
            14'h2fde: oData <= 16'h0000;
            14'h2fdf: oData <= 16'h0000;
            14'h2fe0: oData <= 16'h0000;
            14'h2fe1: oData <= 16'h0000;
            14'h2fe2: oData <= 16'h0000;
            14'h2fe3: oData <= 16'h0000;
            14'h2fe4: oData <= 16'h0000;
            14'h2fe5: oData <= 16'h0000;
            14'h2fe6: oData <= 16'h0000;
            14'h2fe7: oData <= 16'h0000;
            14'h2fe8: oData <= 16'h0000;
            14'h2fe9: oData <= 16'h0000;
            14'h2fea: oData <= 16'h0000;
            14'h2feb: oData <= 16'h0000;
            14'h2fec: oData <= 16'h0000;
            14'h2fed: oData <= 16'h0000;
            14'h2fee: oData <= 16'h0000;
            14'h2fef: oData <= 16'h0000;
            14'h2ff0: oData <= 16'h0000;
            14'h2ff1: oData <= 16'h0000;
            14'h2ff2: oData <= 16'h0000;
            14'h2ff3: oData <= 16'h0000;
            14'h2ff4: oData <= 16'h0000;
            14'h2ff5: oData <= 16'h0000;
            14'h2ff6: oData <= 16'h0000;
            14'h2ff7: oData <= 16'h0000;
            14'h2ff8: oData <= 16'h0000;
            14'h2ff9: oData <= 16'h0000;
            14'h2ffa: oData <= 16'h0000;
            14'h2ffb: oData <= 16'h0000;
            14'h2ffc: oData <= 16'h0000;
            14'h2ffd: oData <= 16'h0000;
            14'h2ffe: oData <= 16'h0000;
            14'h2fff: oData <= 16'h0000;
            14'h3000: oData <= 16'h0000;
            14'h3001: oData <= 16'h0000;
            14'h3002: oData <= 16'h0000;
            14'h3003: oData <= 16'h0000;
            14'h3004: oData <= 16'h0000;
            14'h3005: oData <= 16'h0000;
            14'h3006: oData <= 16'h0000;
            14'h3007: oData <= 16'h0000;
            14'h3008: oData <= 16'h0000;
            14'h3009: oData <= 16'h0000;
            14'h300a: oData <= 16'h0000;
            14'h300b: oData <= 16'h0000;
            14'h300c: oData <= 16'h0000;
            14'h300d: oData <= 16'h0000;
            14'h300e: oData <= 16'h0000;
            14'h300f: oData <= 16'h0000;
            14'h3010: oData <= 16'h0000;
            14'h3011: oData <= 16'h0000;
            14'h3012: oData <= 16'h0000;
            14'h3013: oData <= 16'h0000;
            14'h3014: oData <= 16'h0000;
            14'h3015: oData <= 16'h0000;
            14'h3016: oData <= 16'h0000;
            14'h3017: oData <= 16'h0000;
            14'h3018: oData <= 16'h0000;
            14'h3019: oData <= 16'h0000;
            14'h301a: oData <= 16'h0000;
            14'h301b: oData <= 16'h0000;
            14'h301c: oData <= 16'h0000;
            14'h301d: oData <= 16'h0000;
            14'h301e: oData <= 16'h0000;
            14'h301f: oData <= 16'h0000;
            14'h3020: oData <= 16'h0000;
            14'h3021: oData <= 16'h0000;
            14'h3022: oData <= 16'h0000;
            14'h3023: oData <= 16'h0000;
            14'h3024: oData <= 16'h0000;
            14'h3025: oData <= 16'h0000;
            14'h3026: oData <= 16'h0000;
            14'h3027: oData <= 16'h0000;
            14'h3028: oData <= 16'h0000;
            14'h3029: oData <= 16'h0000;
            14'h302a: oData <= 16'h0000;
            14'h302b: oData <= 16'h0000;
            14'h302c: oData <= 16'h0000;
            14'h302d: oData <= 16'h0000;
            14'h302e: oData <= 16'h0000;
            14'h302f: oData <= 16'h0000;
            14'h3030: oData <= 16'h0000;
            14'h3031: oData <= 16'h0000;
            14'h3032: oData <= 16'h0000;
            14'h3033: oData <= 16'h0000;
            14'h3034: oData <= 16'h0000;
            14'h3035: oData <= 16'h0000;
            14'h3036: oData <= 16'h0000;
            14'h3037: oData <= 16'h0000;
            14'h3038: oData <= 16'h0000;
            14'h3039: oData <= 16'h0000;
            14'h303a: oData <= 16'h0000;
            14'h303b: oData <= 16'h0000;
            14'h303c: oData <= 16'h0000;
            14'h303d: oData <= 16'h0000;
            14'h303e: oData <= 16'h0000;
            14'h303f: oData <= 16'h0000;
            14'h3040: oData <= 16'h0000;
            14'h3041: oData <= 16'h0000;
            14'h3042: oData <= 16'h0000;
            14'h3043: oData <= 16'h0000;
            14'h3044: oData <= 16'h0000;
            14'h3045: oData <= 16'h0000;
            14'h3046: oData <= 16'h0000;
            14'h3047: oData <= 16'h0000;
            14'h3048: oData <= 16'h0000;
            14'h3049: oData <= 16'h0000;
            14'h304a: oData <= 16'h0000;
            14'h304b: oData <= 16'h0000;
            14'h304c: oData <= 16'h0000;
            14'h304d: oData <= 16'h0000;
            14'h304e: oData <= 16'h0000;
            14'h304f: oData <= 16'h0000;
            14'h3050: oData <= 16'h0000;
            14'h3051: oData <= 16'h0000;
            14'h3052: oData <= 16'h0000;
            14'h3053: oData <= 16'h0000;
            14'h3054: oData <= 16'h0000;
            14'h3055: oData <= 16'h0000;
            14'h3056: oData <= 16'h0000;
            14'h3057: oData <= 16'h0000;
            14'h3058: oData <= 16'h0000;
            14'h3059: oData <= 16'h0000;
            14'h305a: oData <= 16'h0000;
            14'h305b: oData <= 16'h0000;
            14'h305c: oData <= 16'h0000;
            14'h305d: oData <= 16'h0000;
            14'h305e: oData <= 16'h0000;
            14'h305f: oData <= 16'h0000;
            14'h3060: oData <= 16'h0000;
            14'h3061: oData <= 16'h0000;
            14'h3062: oData <= 16'h0000;
            14'h3063: oData <= 16'h0000;
            14'h3064: oData <= 16'h0000;
            14'h3065: oData <= 16'h0000;
            14'h3066: oData <= 16'h0000;
            14'h3067: oData <= 16'h0000;
            14'h3068: oData <= 16'h0000;
            14'h3069: oData <= 16'h0000;
            14'h306a: oData <= 16'h0000;
            14'h306b: oData <= 16'h0000;
            14'h306c: oData <= 16'h0000;
            14'h306d: oData <= 16'h0000;
            14'h306e: oData <= 16'h0000;
            14'h306f: oData <= 16'h0000;
            14'h3070: oData <= 16'h0000;
            14'h3071: oData <= 16'h0000;
            14'h3072: oData <= 16'h0000;
            14'h3073: oData <= 16'h0000;
            14'h3074: oData <= 16'h0000;
            14'h3075: oData <= 16'h0000;
            14'h3076: oData <= 16'h0000;
            14'h3077: oData <= 16'h0000;
            14'h3078: oData <= 16'h0000;
            14'h3079: oData <= 16'h0000;
            14'h307a: oData <= 16'h0000;
            14'h307b: oData <= 16'h0000;
            14'h307c: oData <= 16'h0000;
            14'h307d: oData <= 16'h0000;
            14'h307e: oData <= 16'h0000;
            14'h307f: oData <= 16'h0000;
            14'h3080: oData <= 16'h0000;
            14'h3081: oData <= 16'h0000;
            14'h3082: oData <= 16'h0000;
            14'h3083: oData <= 16'h0000;
            14'h3084: oData <= 16'h0000;
            14'h3085: oData <= 16'h0000;
            14'h3086: oData <= 16'h0000;
            14'h3087: oData <= 16'h0000;
            14'h3088: oData <= 16'h0000;
            14'h3089: oData <= 16'h0000;
            14'h308a: oData <= 16'h0000;
            14'h308b: oData <= 16'h0000;
            14'h308c: oData <= 16'h0000;
            14'h308d: oData <= 16'h0000;
            14'h308e: oData <= 16'h0000;
            14'h308f: oData <= 16'h0000;
            14'h3090: oData <= 16'h0000;
            14'h3091: oData <= 16'h0000;
            14'h3092: oData <= 16'h0000;
            14'h3093: oData <= 16'h0000;
            14'h3094: oData <= 16'h0000;
            14'h3095: oData <= 16'h0000;
            14'h3096: oData <= 16'h0000;
            14'h3097: oData <= 16'h0000;
            14'h3098: oData <= 16'h0000;
            14'h3099: oData <= 16'h0000;
            14'h309a: oData <= 16'h0000;
            14'h309b: oData <= 16'h0000;
            14'h309c: oData <= 16'h0000;
            14'h309d: oData <= 16'h0000;
            14'h309e: oData <= 16'h0000;
            14'h309f: oData <= 16'h0000;
            14'h30a0: oData <= 16'h0000;
            14'h30a1: oData <= 16'h0000;
            14'h30a2: oData <= 16'h0000;
            14'h30a3: oData <= 16'h0000;
            14'h30a4: oData <= 16'h0000;
            14'h30a5: oData <= 16'h0000;
            14'h30a6: oData <= 16'h0000;
            14'h30a7: oData <= 16'h0000;
            14'h30a8: oData <= 16'h0000;
            14'h30a9: oData <= 16'h0000;
            14'h30aa: oData <= 16'h0000;
            14'h30ab: oData <= 16'h0000;
            14'h30ac: oData <= 16'h0000;
            14'h30ad: oData <= 16'h0000;
            14'h30ae: oData <= 16'h0000;
            14'h30af: oData <= 16'h0000;
            14'h30b0: oData <= 16'h0000;
            14'h30b1: oData <= 16'h0000;
            14'h30b2: oData <= 16'h0000;
            14'h30b3: oData <= 16'h0000;
            14'h30b4: oData <= 16'h0000;
            14'h30b5: oData <= 16'h0000;
            14'h30b6: oData <= 16'h0000;
            14'h30b7: oData <= 16'h0000;
            14'h30b8: oData <= 16'h0000;
            14'h30b9: oData <= 16'h0000;
            14'h30ba: oData <= 16'h0000;
            14'h30bb: oData <= 16'h0000;
            14'h30bc: oData <= 16'h0000;
            14'h30bd: oData <= 16'h0000;
            14'h30be: oData <= 16'h0000;
            14'h30bf: oData <= 16'h0000;
            14'h30c0: oData <= 16'h0000;
            14'h30c1: oData <= 16'h0000;
            14'h30c2: oData <= 16'h0000;
            14'h30c3: oData <= 16'h0000;
            14'h30c4: oData <= 16'h0000;
            14'h30c5: oData <= 16'h0000;
            14'h30c6: oData <= 16'h0000;
            14'h30c7: oData <= 16'h0000;
            14'h30c8: oData <= 16'h0000;
            14'h30c9: oData <= 16'h0000;
            14'h30ca: oData <= 16'h0000;
            14'h30cb: oData <= 16'h0000;
            14'h30cc: oData <= 16'h0000;
            14'h30cd: oData <= 16'h0000;
            14'h30ce: oData <= 16'h0000;
            14'h30cf: oData <= 16'h0000;
            14'h30d0: oData <= 16'h0000;
            14'h30d1: oData <= 16'h0000;
            14'h30d2: oData <= 16'h0000;
            14'h30d3: oData <= 16'h0000;
            14'h30d4: oData <= 16'h0000;
            14'h30d5: oData <= 16'h0000;
            14'h30d6: oData <= 16'h0000;
            14'h30d7: oData <= 16'h0000;
            14'h30d8: oData <= 16'h0000;
            14'h30d9: oData <= 16'h0000;
            14'h30da: oData <= 16'h0000;
            14'h30db: oData <= 16'h0000;
            14'h30dc: oData <= 16'h0000;
            14'h30dd: oData <= 16'h0000;
            14'h30de: oData <= 16'h0000;
            14'h30df: oData <= 16'h0000;
            14'h30e0: oData <= 16'h0000;
            14'h30e1: oData <= 16'h0000;
            14'h30e2: oData <= 16'h0000;
            14'h30e3: oData <= 16'h0000;
            14'h30e4: oData <= 16'h0000;
            14'h30e5: oData <= 16'h0000;
            14'h30e6: oData <= 16'h0000;
            14'h30e7: oData <= 16'h0000;
            14'h30e8: oData <= 16'h0000;
            14'h30e9: oData <= 16'h0000;
            14'h30ea: oData <= 16'h0000;
            14'h30eb: oData <= 16'h0000;
            14'h30ec: oData <= 16'h0000;
            14'h30ed: oData <= 16'h0000;
            14'h30ee: oData <= 16'h0000;
            14'h30ef: oData <= 16'h0000;
            14'h30f0: oData <= 16'h0000;
            14'h30f1: oData <= 16'h0000;
            14'h30f2: oData <= 16'h0000;
            14'h30f3: oData <= 16'h0000;
            14'h30f4: oData <= 16'h0000;
            14'h30f5: oData <= 16'h0000;
            14'h30f6: oData <= 16'h0000;
            14'h30f7: oData <= 16'h0000;
            14'h30f8: oData <= 16'h0000;
            14'h30f9: oData <= 16'h0000;
            14'h30fa: oData <= 16'h0000;
            14'h30fb: oData <= 16'h0000;
            14'h30fc: oData <= 16'h0000;
            14'h30fd: oData <= 16'h0000;
            14'h30fe: oData <= 16'h0000;
            14'h30ff: oData <= 16'h0000;
            14'h3100: oData <= 16'h0000;
            14'h3101: oData <= 16'h0000;
            14'h3102: oData <= 16'h0000;
            14'h3103: oData <= 16'h0000;
            14'h3104: oData <= 16'h0000;
            14'h3105: oData <= 16'h0000;
            14'h3106: oData <= 16'h0000;
            14'h3107: oData <= 16'h0000;
            14'h3108: oData <= 16'h0000;
            14'h3109: oData <= 16'h0000;
            14'h310a: oData <= 16'h0000;
            14'h310b: oData <= 16'h0000;
            14'h310c: oData <= 16'h0000;
            14'h310d: oData <= 16'h0000;
            14'h310e: oData <= 16'h0000;
            14'h310f: oData <= 16'h0000;
            14'h3110: oData <= 16'h0000;
            14'h3111: oData <= 16'h0000;
            14'h3112: oData <= 16'h0000;
            14'h3113: oData <= 16'h0000;
            14'h3114: oData <= 16'h0000;
            14'h3115: oData <= 16'h0000;
            14'h3116: oData <= 16'h0000;
            14'h3117: oData <= 16'h0000;
            14'h3118: oData <= 16'h0000;
            14'h3119: oData <= 16'h0000;
            14'h311a: oData <= 16'h0000;
            14'h311b: oData <= 16'h0000;
            14'h311c: oData <= 16'h0000;
            14'h311d: oData <= 16'h0000;
            14'h311e: oData <= 16'h0000;
            14'h311f: oData <= 16'h0000;
            14'h3120: oData <= 16'h0000;
            14'h3121: oData <= 16'h0000;
            14'h3122: oData <= 16'h0000;
            14'h3123: oData <= 16'h0000;
            14'h3124: oData <= 16'h0000;
            14'h3125: oData <= 16'h0000;
            14'h3126: oData <= 16'h0000;
            14'h3127: oData <= 16'h0000;
            14'h3128: oData <= 16'h0000;
            14'h3129: oData <= 16'h0000;
            14'h312a: oData <= 16'h0000;
            14'h312b: oData <= 16'h0000;
            14'h312c: oData <= 16'h0000;
            14'h312d: oData <= 16'h0000;
            14'h312e: oData <= 16'h0000;
            14'h312f: oData <= 16'h0000;
            14'h3130: oData <= 16'h0000;
            14'h3131: oData <= 16'h0000;
            14'h3132: oData <= 16'h0000;
            14'h3133: oData <= 16'h0000;
            14'h3134: oData <= 16'h0000;
            14'h3135: oData <= 16'h0000;
            14'h3136: oData <= 16'h0000;
            14'h3137: oData <= 16'h0000;
            14'h3138: oData <= 16'h0000;
            14'h3139: oData <= 16'h0000;
            14'h313a: oData <= 16'h0000;
            14'h313b: oData <= 16'h0000;
            14'h313c: oData <= 16'h0000;
            14'h313d: oData <= 16'h0000;
            14'h313e: oData <= 16'h0000;
            14'h313f: oData <= 16'h0000;
            14'h3140: oData <= 16'h0000;
            14'h3141: oData <= 16'h0000;
            14'h3142: oData <= 16'h0000;
            14'h3143: oData <= 16'h0000;
            14'h3144: oData <= 16'h0000;
            14'h3145: oData <= 16'h0000;
            14'h3146: oData <= 16'h0000;
            14'h3147: oData <= 16'h0000;
            14'h3148: oData <= 16'h0000;
            14'h3149: oData <= 16'h0000;
            14'h314a: oData <= 16'h0000;
            14'h314b: oData <= 16'h0000;
            14'h314c: oData <= 16'h0000;
            14'h314d: oData <= 16'h0000;
            14'h314e: oData <= 16'h0000;
            14'h314f: oData <= 16'h0000;
            14'h3150: oData <= 16'h0000;
            14'h3151: oData <= 16'h0000;
            14'h3152: oData <= 16'h0000;
            14'h3153: oData <= 16'h0000;
            14'h3154: oData <= 16'h0000;
            14'h3155: oData <= 16'h0000;
            14'h3156: oData <= 16'h0000;
            14'h3157: oData <= 16'h0000;
            14'h3158: oData <= 16'h0000;
            14'h3159: oData <= 16'h0000;
            14'h315a: oData <= 16'h0000;
            14'h315b: oData <= 16'h0000;
            14'h315c: oData <= 16'h0000;
            14'h315d: oData <= 16'h0000;
            14'h315e: oData <= 16'h0000;
            14'h315f: oData <= 16'h0000;
            14'h3160: oData <= 16'h0000;
            14'h3161: oData <= 16'h0000;
            14'h3162: oData <= 16'h0000;
            14'h3163: oData <= 16'h0000;
            14'h3164: oData <= 16'h0000;
            14'h3165: oData <= 16'h0000;
            14'h3166: oData <= 16'h0000;
            14'h3167: oData <= 16'h0000;
            14'h3168: oData <= 16'h0000;
            14'h3169: oData <= 16'h0000;
            14'h316a: oData <= 16'h0000;
            14'h316b: oData <= 16'h0000;
            14'h316c: oData <= 16'h0000;
            14'h316d: oData <= 16'h0000;
            14'h316e: oData <= 16'h0000;
            14'h316f: oData <= 16'h0000;
            14'h3170: oData <= 16'h0000;
            14'h3171: oData <= 16'h0000;
            14'h3172: oData <= 16'h0000;
            14'h3173: oData <= 16'h0000;
            14'h3174: oData <= 16'h0000;
            14'h3175: oData <= 16'h0000;
            14'h3176: oData <= 16'h0000;
            14'h3177: oData <= 16'h0000;
            14'h3178: oData <= 16'h0000;
            14'h3179: oData <= 16'h0000;
            14'h317a: oData <= 16'h0000;
            14'h317b: oData <= 16'h0000;
            14'h317c: oData <= 16'h0000;
            14'h317d: oData <= 16'h0000;
            14'h317e: oData <= 16'h0000;
            14'h317f: oData <= 16'h0000;
            14'h3180: oData <= 16'h0000;
            14'h3181: oData <= 16'h0000;
            14'h3182: oData <= 16'h0000;
            14'h3183: oData <= 16'h0000;
            14'h3184: oData <= 16'h0000;
            14'h3185: oData <= 16'h0000;
            14'h3186: oData <= 16'h0000;
            14'h3187: oData <= 16'h0000;
            14'h3188: oData <= 16'h0000;
            14'h3189: oData <= 16'h0000;
            14'h318a: oData <= 16'h0000;
            14'h318b: oData <= 16'h0000;
            14'h318c: oData <= 16'h0000;
            14'h318d: oData <= 16'h0000;
            14'h318e: oData <= 16'h0000;
            14'h318f: oData <= 16'h0000;
            14'h3190: oData <= 16'h0000;
            14'h3191: oData <= 16'h0000;
            14'h3192: oData <= 16'h0000;
            14'h3193: oData <= 16'h0000;
            14'h3194: oData <= 16'h0000;
            14'h3195: oData <= 16'h0000;
            14'h3196: oData <= 16'h0000;
            14'h3197: oData <= 16'h0000;
            14'h3198: oData <= 16'h0000;
            14'h3199: oData <= 16'h0000;
            14'h319a: oData <= 16'h0000;
            14'h319b: oData <= 16'h0000;
            14'h319c: oData <= 16'h0000;
            14'h319d: oData <= 16'h0000;
            14'h319e: oData <= 16'h0000;
            14'h319f: oData <= 16'h0000;
            14'h31a0: oData <= 16'h0000;
            14'h31a1: oData <= 16'h0000;
            14'h31a2: oData <= 16'h0000;
            14'h31a3: oData <= 16'h0000;
            14'h31a4: oData <= 16'h0000;
            14'h31a5: oData <= 16'h0000;
            14'h31a6: oData <= 16'h0000;
            14'h31a7: oData <= 16'h0000;
            14'h31a8: oData <= 16'h0000;
            14'h31a9: oData <= 16'h0000;
            14'h31aa: oData <= 16'h0000;
            14'h31ab: oData <= 16'h0000;
            14'h31ac: oData <= 16'h0000;
            14'h31ad: oData <= 16'h0000;
            14'h31ae: oData <= 16'h0000;
            14'h31af: oData <= 16'h0000;
            14'h31b0: oData <= 16'h0000;
            14'h31b1: oData <= 16'h0000;
            14'h31b2: oData <= 16'h0000;
            14'h31b3: oData <= 16'h0000;
            14'h31b4: oData <= 16'h0000;
            14'h31b5: oData <= 16'h0000;
            14'h31b6: oData <= 16'h0000;
            14'h31b7: oData <= 16'h0000;
            14'h31b8: oData <= 16'h0000;
            14'h31b9: oData <= 16'h0000;
            14'h31ba: oData <= 16'h0000;
            14'h31bb: oData <= 16'h0000;
            14'h31bc: oData <= 16'h0000;
            14'h31bd: oData <= 16'h0000;
            14'h31be: oData <= 16'h0000;
            14'h31bf: oData <= 16'h0000;
            14'h31c0: oData <= 16'h0000;
            14'h31c1: oData <= 16'h0000;
            14'h31c2: oData <= 16'h0000;
            14'h31c3: oData <= 16'h0000;
            14'h31c4: oData <= 16'h0000;
            14'h31c5: oData <= 16'h0000;
            14'h31c6: oData <= 16'h0000;
            14'h31c7: oData <= 16'h0000;
            14'h31c8: oData <= 16'h0000;
            14'h31c9: oData <= 16'h0000;
            14'h31ca: oData <= 16'h0000;
            14'h31cb: oData <= 16'h0000;
            14'h31cc: oData <= 16'h0000;
            14'h31cd: oData <= 16'h0000;
            14'h31ce: oData <= 16'h0000;
            14'h31cf: oData <= 16'h0000;
            14'h31d0: oData <= 16'h0000;
            14'h31d1: oData <= 16'h0000;
            14'h31d2: oData <= 16'h0000;
            14'h31d3: oData <= 16'h0000;
            14'h31d4: oData <= 16'h0000;
            14'h31d5: oData <= 16'h0000;
            14'h31d6: oData <= 16'h0000;
            14'h31d7: oData <= 16'h0000;
            14'h31d8: oData <= 16'h0000;
            14'h31d9: oData <= 16'h0000;
            14'h31da: oData <= 16'h0000;
            14'h31db: oData <= 16'h0000;
            14'h31dc: oData <= 16'h0000;
            14'h31dd: oData <= 16'h0000;
            14'h31de: oData <= 16'h0000;
            14'h31df: oData <= 16'h0000;
            14'h31e0: oData <= 16'h0000;
            14'h31e1: oData <= 16'h0000;
            14'h31e2: oData <= 16'h0000;
            14'h31e3: oData <= 16'h0000;
            14'h31e4: oData <= 16'h0000;
            14'h31e5: oData <= 16'h0000;
            14'h31e6: oData <= 16'h0000;
            14'h31e7: oData <= 16'h0000;
            14'h31e8: oData <= 16'h0000;
            14'h31e9: oData <= 16'h0000;
            14'h31ea: oData <= 16'h0000;
            14'h31eb: oData <= 16'h0000;
            14'h31ec: oData <= 16'h0000;
            14'h31ed: oData <= 16'h0000;
            14'h31ee: oData <= 16'h0000;
            14'h31ef: oData <= 16'h0000;
            14'h31f0: oData <= 16'h0000;
            14'h31f1: oData <= 16'h0000;
            14'h31f2: oData <= 16'h0000;
            14'h31f3: oData <= 16'h0000;
            14'h31f4: oData <= 16'h0000;
            14'h31f5: oData <= 16'h0000;
            14'h31f6: oData <= 16'h0000;
            14'h31f7: oData <= 16'h0000;
            14'h31f8: oData <= 16'h0000;
            14'h31f9: oData <= 16'h0000;
            14'h31fa: oData <= 16'h0000;
            14'h31fb: oData <= 16'h0000;
            14'h31fc: oData <= 16'h0000;
            14'h31fd: oData <= 16'h0000;
            14'h31fe: oData <= 16'h0000;
            14'h31ff: oData <= 16'h0000;
            14'h3200: oData <= 16'h0000;
            14'h3201: oData <= 16'h0000;
            14'h3202: oData <= 16'h0000;
            14'h3203: oData <= 16'h0000;
            14'h3204: oData <= 16'h0000;
            14'h3205: oData <= 16'h0000;
            14'h3206: oData <= 16'h0000;
            14'h3207: oData <= 16'h0000;
            14'h3208: oData <= 16'h0000;
            14'h3209: oData <= 16'h0000;
            14'h320a: oData <= 16'h0000;
            14'h320b: oData <= 16'h0000;
            14'h320c: oData <= 16'h0000;
            14'h320d: oData <= 16'h0000;
            14'h320e: oData <= 16'h0000;
            14'h320f: oData <= 16'h0000;
            14'h3210: oData <= 16'h0000;
            14'h3211: oData <= 16'h0000;
            14'h3212: oData <= 16'h0000;
            14'h3213: oData <= 16'h0000;
            14'h3214: oData <= 16'h0000;
            14'h3215: oData <= 16'h0000;
            14'h3216: oData <= 16'h0000;
            14'h3217: oData <= 16'h0000;
            14'h3218: oData <= 16'h0000;
            14'h3219: oData <= 16'h0000;
            14'h321a: oData <= 16'h0000;
            14'h321b: oData <= 16'h0000;
            14'h321c: oData <= 16'h0000;
            14'h321d: oData <= 16'h0000;
            14'h321e: oData <= 16'h0000;
            14'h321f: oData <= 16'h0000;
            14'h3220: oData <= 16'h0000;
            14'h3221: oData <= 16'h0000;
            14'h3222: oData <= 16'h0000;
            14'h3223: oData <= 16'h0000;
            14'h3224: oData <= 16'h0000;
            14'h3225: oData <= 16'h0000;
            14'h3226: oData <= 16'h0000;
            14'h3227: oData <= 16'h0000;
            14'h3228: oData <= 16'h0000;
            14'h3229: oData <= 16'h0000;
            14'h322a: oData <= 16'h0000;
            14'h322b: oData <= 16'h0000;
            14'h322c: oData <= 16'h0000;
            14'h322d: oData <= 16'h0000;
            14'h322e: oData <= 16'h0000;
            14'h322f: oData <= 16'h0000;
            14'h3230: oData <= 16'h0000;
            14'h3231: oData <= 16'h0000;
            14'h3232: oData <= 16'h0000;
            14'h3233: oData <= 16'h0000;
            14'h3234: oData <= 16'h0000;
            14'h3235: oData <= 16'h0000;
            14'h3236: oData <= 16'h0000;
            14'h3237: oData <= 16'h0000;
            14'h3238: oData <= 16'h0000;
            14'h3239: oData <= 16'h0000;
            14'h323a: oData <= 16'h0000;
            14'h323b: oData <= 16'h0000;
            14'h323c: oData <= 16'h0000;
            14'h323d: oData <= 16'h0000;
            14'h323e: oData <= 16'h0000;
            14'h323f: oData <= 16'h0000;
            14'h3240: oData <= 16'h0000;
            14'h3241: oData <= 16'h0000;
            14'h3242: oData <= 16'h0000;
            14'h3243: oData <= 16'h0000;
            14'h3244: oData <= 16'h0000;
            14'h3245: oData <= 16'h0000;
            14'h3246: oData <= 16'h0000;
            14'h3247: oData <= 16'h0000;
            14'h3248: oData <= 16'h0000;
            14'h3249: oData <= 16'h0000;
            14'h324a: oData <= 16'h0000;
            14'h324b: oData <= 16'h0000;
            14'h324c: oData <= 16'h0000;
            14'h324d: oData <= 16'h0000;
            14'h324e: oData <= 16'h0000;
            14'h324f: oData <= 16'h0000;
            14'h3250: oData <= 16'h0000;
            14'h3251: oData <= 16'h0000;
            14'h3252: oData <= 16'h0000;
            14'h3253: oData <= 16'h0000;
            14'h3254: oData <= 16'h0000;
            14'h3255: oData <= 16'h0000;
            14'h3256: oData <= 16'h0000;
            14'h3257: oData <= 16'h0000;
            14'h3258: oData <= 16'h0000;
            14'h3259: oData <= 16'h0000;
            14'h325a: oData <= 16'h0000;
            14'h325b: oData <= 16'h0000;
            14'h325c: oData <= 16'h0000;
            14'h325d: oData <= 16'h0000;
            14'h325e: oData <= 16'h0000;
            14'h325f: oData <= 16'h0000;
            14'h3260: oData <= 16'h0000;
            14'h3261: oData <= 16'h0000;
            14'h3262: oData <= 16'h0000;
            14'h3263: oData <= 16'h0000;
            14'h3264: oData <= 16'h0000;
            14'h3265: oData <= 16'h0000;
            14'h3266: oData <= 16'h0000;
            14'h3267: oData <= 16'h0000;
            14'h3268: oData <= 16'h0000;
            14'h3269: oData <= 16'h0000;
            14'h326a: oData <= 16'h0000;
            14'h326b: oData <= 16'h0000;
            14'h326c: oData <= 16'h0000;
            14'h326d: oData <= 16'h0000;
            14'h326e: oData <= 16'h0000;
            14'h326f: oData <= 16'h0000;
            14'h3270: oData <= 16'h0000;
            14'h3271: oData <= 16'h0000;
            14'h3272: oData <= 16'h0000;
            14'h3273: oData <= 16'h0000;
            14'h3274: oData <= 16'h0000;
            14'h3275: oData <= 16'h0000;
            14'h3276: oData <= 16'h0000;
            14'h3277: oData <= 16'h0000;
            14'h3278: oData <= 16'h0000;
            14'h3279: oData <= 16'h0000;
            14'h327a: oData <= 16'h0000;
            14'h327b: oData <= 16'h0000;
            14'h327c: oData <= 16'h0000;
            14'h327d: oData <= 16'h0000;
            14'h327e: oData <= 16'h0000;
            14'h327f: oData <= 16'h0000;
            14'h3280: oData <= 16'h0000;
            14'h3281: oData <= 16'h0000;
            14'h3282: oData <= 16'h0000;
            14'h3283: oData <= 16'h0000;
            14'h3284: oData <= 16'h0000;
            14'h3285: oData <= 16'h0000;
            14'h3286: oData <= 16'h0000;
            14'h3287: oData <= 16'h0000;
            14'h3288: oData <= 16'h0000;
            14'h3289: oData <= 16'h0000;
            14'h328a: oData <= 16'h0000;
            14'h328b: oData <= 16'h0000;
            14'h328c: oData <= 16'h0000;
            14'h328d: oData <= 16'h0000;
            14'h328e: oData <= 16'h0000;
            14'h328f: oData <= 16'h0000;
            14'h3290: oData <= 16'h0000;
            14'h3291: oData <= 16'h0000;
            14'h3292: oData <= 16'h0000;
            14'h3293: oData <= 16'h0000;
            14'h3294: oData <= 16'h0000;
            14'h3295: oData <= 16'h0000;
            14'h3296: oData <= 16'h0000;
            14'h3297: oData <= 16'h0000;
            14'h3298: oData <= 16'h0000;
            14'h3299: oData <= 16'h0000;
            14'h329a: oData <= 16'h0000;
            14'h329b: oData <= 16'h0000;
            14'h329c: oData <= 16'h0000;
            14'h329d: oData <= 16'h0000;
            14'h329e: oData <= 16'h0000;
            14'h329f: oData <= 16'h0000;
            14'h32a0: oData <= 16'h0000;
            14'h32a1: oData <= 16'h0000;
            14'h32a2: oData <= 16'h0000;
            14'h32a3: oData <= 16'h0000;
            14'h32a4: oData <= 16'h0000;
            14'h32a5: oData <= 16'h0000;
            14'h32a6: oData <= 16'h0000;
            14'h32a7: oData <= 16'h0000;
            14'h32a8: oData <= 16'h0000;
            14'h32a9: oData <= 16'h0000;
            14'h32aa: oData <= 16'h0000;
            14'h32ab: oData <= 16'h0000;
            14'h32ac: oData <= 16'h0000;
            14'h32ad: oData <= 16'h0000;
            14'h32ae: oData <= 16'h0000;
            14'h32af: oData <= 16'h0000;
            14'h32b0: oData <= 16'h0000;
            14'h32b1: oData <= 16'h0000;
            14'h32b2: oData <= 16'h0000;
            14'h32b3: oData <= 16'h0000;
            14'h32b4: oData <= 16'h0000;
            14'h32b5: oData <= 16'h0000;
            14'h32b6: oData <= 16'h0000;
            14'h32b7: oData <= 16'h0000;
            14'h32b8: oData <= 16'h0000;
            14'h32b9: oData <= 16'h0000;
            14'h32ba: oData <= 16'h0000;
            14'h32bb: oData <= 16'h0000;
            14'h32bc: oData <= 16'h0000;
            14'h32bd: oData <= 16'h0000;
            14'h32be: oData <= 16'h0000;
            14'h32bf: oData <= 16'h0000;
            14'h32c0: oData <= 16'h0000;
            14'h32c1: oData <= 16'h0000;
            14'h32c2: oData <= 16'h0000;
            14'h32c3: oData <= 16'h0000;
            14'h32c4: oData <= 16'h0000;
            14'h32c5: oData <= 16'h0000;
            14'h32c6: oData <= 16'h0000;
            14'h32c7: oData <= 16'h0000;
            14'h32c8: oData <= 16'h0000;
            14'h32c9: oData <= 16'h0000;
            14'h32ca: oData <= 16'h0000;
            14'h32cb: oData <= 16'h0000;
            14'h32cc: oData <= 16'h0000;
            14'h32cd: oData <= 16'h0000;
            14'h32ce: oData <= 16'h0000;
            14'h32cf: oData <= 16'h0000;
            14'h32d0: oData <= 16'h0000;
            14'h32d1: oData <= 16'h0000;
            14'h32d2: oData <= 16'h0000;
            14'h32d3: oData <= 16'h0000;
            14'h32d4: oData <= 16'h0000;
            14'h32d5: oData <= 16'h0000;
            14'h32d6: oData <= 16'h0000;
            14'h32d7: oData <= 16'h0000;
            14'h32d8: oData <= 16'h0000;
            14'h32d9: oData <= 16'h0000;
            14'h32da: oData <= 16'h0000;
            14'h32db: oData <= 16'h0000;
            14'h32dc: oData <= 16'h0000;
            14'h32dd: oData <= 16'h0000;
            14'h32de: oData <= 16'h0000;
            14'h32df: oData <= 16'h0000;
            14'h32e0: oData <= 16'h0000;
            14'h32e1: oData <= 16'h0000;
            14'h32e2: oData <= 16'h0000;
            14'h32e3: oData <= 16'h0000;
            14'h32e4: oData <= 16'h0000;
            14'h32e5: oData <= 16'h0000;
            14'h32e6: oData <= 16'h0000;
            14'h32e7: oData <= 16'h0000;
            14'h32e8: oData <= 16'h0000;
            14'h32e9: oData <= 16'h0000;
            14'h32ea: oData <= 16'h0000;
            14'h32eb: oData <= 16'h0000;
            14'h32ec: oData <= 16'h0000;
            14'h32ed: oData <= 16'h0000;
            14'h32ee: oData <= 16'h0000;
            14'h32ef: oData <= 16'h0000;
            14'h32f0: oData <= 16'h0000;
            14'h32f1: oData <= 16'h0000;
            14'h32f2: oData <= 16'h0000;
            14'h32f3: oData <= 16'h0000;
            14'h32f4: oData <= 16'h0000;
            14'h32f5: oData <= 16'h0000;
            14'h32f6: oData <= 16'h0000;
            14'h32f7: oData <= 16'h0000;
            14'h32f8: oData <= 16'h0000;
            14'h32f9: oData <= 16'h0000;
            14'h32fa: oData <= 16'h0000;
            14'h32fb: oData <= 16'h0000;
            14'h32fc: oData <= 16'h0000;
            14'h32fd: oData <= 16'h0000;
            14'h32fe: oData <= 16'h0000;
            14'h32ff: oData <= 16'h0000;
            14'h3300: oData <= 16'h0000;
            14'h3301: oData <= 16'h0000;
            14'h3302: oData <= 16'h0000;
            14'h3303: oData <= 16'h0000;
            14'h3304: oData <= 16'h0000;
            14'h3305: oData <= 16'h0000;
            14'h3306: oData <= 16'h0000;
            14'h3307: oData <= 16'h0000;
            14'h3308: oData <= 16'h0000;
            14'h3309: oData <= 16'h0000;
            14'h330a: oData <= 16'h0000;
            14'h330b: oData <= 16'h0000;
            14'h330c: oData <= 16'h0000;
            14'h330d: oData <= 16'h0000;
            14'h330e: oData <= 16'h0000;
            14'h330f: oData <= 16'h0000;
            14'h3310: oData <= 16'h0000;
            14'h3311: oData <= 16'h0000;
            14'h3312: oData <= 16'h0000;
            14'h3313: oData <= 16'h0000;
            14'h3314: oData <= 16'h0000;
            14'h3315: oData <= 16'h0000;
            14'h3316: oData <= 16'h0000;
            14'h3317: oData <= 16'h0000;
            14'h3318: oData <= 16'h0000;
            14'h3319: oData <= 16'h0000;
            14'h331a: oData <= 16'h0000;
            14'h331b: oData <= 16'h0000;
            14'h331c: oData <= 16'h0000;
            14'h331d: oData <= 16'h0000;
            14'h331e: oData <= 16'h0000;
            14'h331f: oData <= 16'h0000;
            14'h3320: oData <= 16'h0000;
            14'h3321: oData <= 16'h0000;
            14'h3322: oData <= 16'h0000;
            14'h3323: oData <= 16'h0000;
            14'h3324: oData <= 16'h0000;
            14'h3325: oData <= 16'h0000;
            14'h3326: oData <= 16'h0000;
            14'h3327: oData <= 16'h0000;
            14'h3328: oData <= 16'h0000;
            14'h3329: oData <= 16'h0000;
            14'h332a: oData <= 16'h0000;
            14'h332b: oData <= 16'h0000;
            14'h332c: oData <= 16'h0000;
            14'h332d: oData <= 16'h0000;
            14'h332e: oData <= 16'h0000;
            14'h332f: oData <= 16'h0000;
            14'h3330: oData <= 16'h0000;
            14'h3331: oData <= 16'h0000;
            14'h3332: oData <= 16'h0000;
            14'h3333: oData <= 16'h0000;
            14'h3334: oData <= 16'h0000;
            14'h3335: oData <= 16'h0000;
            14'h3336: oData <= 16'h0000;
            14'h3337: oData <= 16'h0000;
            14'h3338: oData <= 16'h0000;
            14'h3339: oData <= 16'h0000;
            14'h333a: oData <= 16'h0000;
            14'h333b: oData <= 16'h0000;
            14'h333c: oData <= 16'h0000;
            14'h333d: oData <= 16'h0000;
            14'h333e: oData <= 16'h0000;
            14'h333f: oData <= 16'h0000;
            14'h3340: oData <= 16'h0000;
            14'h3341: oData <= 16'h0000;
            14'h3342: oData <= 16'h0000;
            14'h3343: oData <= 16'h0000;
            14'h3344: oData <= 16'h0000;
            14'h3345: oData <= 16'h0000;
            14'h3346: oData <= 16'h0000;
            14'h3347: oData <= 16'h0000;
            14'h3348: oData <= 16'h0000;
            14'h3349: oData <= 16'h0000;
            14'h334a: oData <= 16'h0000;
            14'h334b: oData <= 16'h0000;
            14'h334c: oData <= 16'h0000;
            14'h334d: oData <= 16'h0000;
            14'h334e: oData <= 16'h0000;
            14'h334f: oData <= 16'h0000;
            14'h3350: oData <= 16'h0000;
            14'h3351: oData <= 16'h0000;
            14'h3352: oData <= 16'h0000;
            14'h3353: oData <= 16'h0000;
            14'h3354: oData <= 16'h0000;
            14'h3355: oData <= 16'h0000;
            14'h3356: oData <= 16'h0000;
            14'h3357: oData <= 16'h0000;
            14'h3358: oData <= 16'h0000;
            14'h3359: oData <= 16'h0000;
            14'h335a: oData <= 16'h0000;
            14'h335b: oData <= 16'h0000;
            14'h335c: oData <= 16'h0000;
            14'h335d: oData <= 16'h0000;
            14'h335e: oData <= 16'h0000;
            14'h335f: oData <= 16'h0000;
            14'h3360: oData <= 16'h0000;
            14'h3361: oData <= 16'h0000;
            14'h3362: oData <= 16'h0000;
            14'h3363: oData <= 16'h0000;
            14'h3364: oData <= 16'h0000;
            14'h3365: oData <= 16'h0000;
            14'h3366: oData <= 16'h0000;
            14'h3367: oData <= 16'h0000;
            14'h3368: oData <= 16'h0000;
            14'h3369: oData <= 16'h0000;
            14'h336a: oData <= 16'h0000;
            14'h336b: oData <= 16'h0000;
            14'h336c: oData <= 16'h0000;
            14'h336d: oData <= 16'h0000;
            14'h336e: oData <= 16'h0000;
            14'h336f: oData <= 16'h0000;
            14'h3370: oData <= 16'h0000;
            14'h3371: oData <= 16'h0000;
            14'h3372: oData <= 16'h0000;
            14'h3373: oData <= 16'h0000;
            14'h3374: oData <= 16'h0000;
            14'h3375: oData <= 16'h0000;
            14'h3376: oData <= 16'h0000;
            14'h3377: oData <= 16'h0000;
            14'h3378: oData <= 16'h0000;
            14'h3379: oData <= 16'h0000;
            14'h337a: oData <= 16'h0000;
            14'h337b: oData <= 16'h0000;
            14'h337c: oData <= 16'h0000;
            14'h337d: oData <= 16'h0000;
            14'h337e: oData <= 16'h0000;
            14'h337f: oData <= 16'h0000;
            14'h3380: oData <= 16'h0000;
            14'h3381: oData <= 16'h0000;
            14'h3382: oData <= 16'h0000;
            14'h3383: oData <= 16'h0000;
            14'h3384: oData <= 16'h0000;
            14'h3385: oData <= 16'h0000;
            14'h3386: oData <= 16'h0000;
            14'h3387: oData <= 16'h0000;
            14'h3388: oData <= 16'h0000;
            14'h3389: oData <= 16'h0000;
            14'h338a: oData <= 16'h0000;
            14'h338b: oData <= 16'h0000;
            14'h338c: oData <= 16'h0000;
            14'h338d: oData <= 16'h0000;
            14'h338e: oData <= 16'h0000;
            14'h338f: oData <= 16'h0000;
            14'h3390: oData <= 16'h0000;
            14'h3391: oData <= 16'h0000;
            14'h3392: oData <= 16'h0000;
            14'h3393: oData <= 16'h0000;
            14'h3394: oData <= 16'h0000;
            14'h3395: oData <= 16'h0000;
            14'h3396: oData <= 16'h0000;
            14'h3397: oData <= 16'h0000;
            14'h3398: oData <= 16'h0000;
            14'h3399: oData <= 16'h0000;
            14'h339a: oData <= 16'h0000;
            14'h339b: oData <= 16'h0000;
            14'h339c: oData <= 16'h0000;
            14'h339d: oData <= 16'h0000;
            14'h339e: oData <= 16'h0000;
            14'h339f: oData <= 16'h0000;
            14'h33a0: oData <= 16'h0000;
            14'h33a1: oData <= 16'h0000;
            14'h33a2: oData <= 16'h0000;
            14'h33a3: oData <= 16'h0000;
            14'h33a4: oData <= 16'h0000;
            14'h33a5: oData <= 16'h0000;
            14'h33a6: oData <= 16'h0000;
            14'h33a7: oData <= 16'h0000;
            14'h33a8: oData <= 16'h0000;
            14'h33a9: oData <= 16'h0000;
            14'h33aa: oData <= 16'h0000;
            14'h33ab: oData <= 16'h0000;
            14'h33ac: oData <= 16'h0000;
            14'h33ad: oData <= 16'h0000;
            14'h33ae: oData <= 16'h0000;
            14'h33af: oData <= 16'h0000;
            14'h33b0: oData <= 16'h0000;
            14'h33b1: oData <= 16'h0000;
            14'h33b2: oData <= 16'h0000;
            14'h33b3: oData <= 16'h0000;
            14'h33b4: oData <= 16'h0000;
            14'h33b5: oData <= 16'h0000;
            14'h33b6: oData <= 16'h0000;
            14'h33b7: oData <= 16'h0000;
            14'h33b8: oData <= 16'h0000;
            14'h33b9: oData <= 16'h0000;
            14'h33ba: oData <= 16'h0000;
            14'h33bb: oData <= 16'h0000;
            14'h33bc: oData <= 16'h0000;
            14'h33bd: oData <= 16'h0000;
            14'h33be: oData <= 16'h0000;
            14'h33bf: oData <= 16'h0000;
            14'h33c0: oData <= 16'h0000;
            14'h33c1: oData <= 16'h0000;
            14'h33c2: oData <= 16'h0000;
            14'h33c3: oData <= 16'h0000;
            14'h33c4: oData <= 16'h0000;
            14'h33c5: oData <= 16'h0000;
            14'h33c6: oData <= 16'h0000;
            14'h33c7: oData <= 16'h0000;
            14'h33c8: oData <= 16'h0000;
            14'h33c9: oData <= 16'h0000;
            14'h33ca: oData <= 16'h0000;
            14'h33cb: oData <= 16'h0000;
            14'h33cc: oData <= 16'h0000;
            14'h33cd: oData <= 16'h0000;
            14'h33ce: oData <= 16'h0000;
            14'h33cf: oData <= 16'h0000;
            14'h33d0: oData <= 16'h0000;
            14'h33d1: oData <= 16'h0000;
            14'h33d2: oData <= 16'h0000;
            14'h33d3: oData <= 16'h0000;
            14'h33d4: oData <= 16'h0000;
            14'h33d5: oData <= 16'h0000;
            14'h33d6: oData <= 16'h0000;
            14'h33d7: oData <= 16'h0000;
            14'h33d8: oData <= 16'h0000;
            14'h33d9: oData <= 16'h0000;
            14'h33da: oData <= 16'h0000;
            14'h33db: oData <= 16'h0000;
            14'h33dc: oData <= 16'h0000;
            14'h33dd: oData <= 16'h0000;
            14'h33de: oData <= 16'h0000;
            14'h33df: oData <= 16'h0000;
            14'h33e0: oData <= 16'h0000;
            14'h33e1: oData <= 16'h0000;
            14'h33e2: oData <= 16'h0000;
            14'h33e3: oData <= 16'h0000;
            14'h33e4: oData <= 16'h0000;
            14'h33e5: oData <= 16'h0000;
            14'h33e6: oData <= 16'h0000;
            14'h33e7: oData <= 16'h0000;
            14'h33e8: oData <= 16'h0000;
            14'h33e9: oData <= 16'h0000;
            14'h33ea: oData <= 16'h0000;
            14'h33eb: oData <= 16'h0000;
            14'h33ec: oData <= 16'h0000;
            14'h33ed: oData <= 16'h0000;
            14'h33ee: oData <= 16'h0000;
            14'h33ef: oData <= 16'h0000;
            14'h33f0: oData <= 16'h0000;
            14'h33f1: oData <= 16'h0000;
            14'h33f2: oData <= 16'h0000;
            14'h33f3: oData <= 16'h0000;
            14'h33f4: oData <= 16'h0000;
            14'h33f5: oData <= 16'h0000;
            14'h33f6: oData <= 16'h0000;
            14'h33f7: oData <= 16'h0000;
            14'h33f8: oData <= 16'h0000;
            14'h33f9: oData <= 16'h0000;
            14'h33fa: oData <= 16'h0000;
            14'h33fb: oData <= 16'h0000;
            14'h33fc: oData <= 16'h0000;
            14'h33fd: oData <= 16'h0000;
            14'h33fe: oData <= 16'h0000;
            14'h33ff: oData <= 16'h0000;
            14'h3400: oData <= 16'h0000;
            14'h3401: oData <= 16'h0000;
            14'h3402: oData <= 16'h0000;
            14'h3403: oData <= 16'h0000;
            14'h3404: oData <= 16'h0000;
            14'h3405: oData <= 16'h0000;
            14'h3406: oData <= 16'h0000;
            14'h3407: oData <= 16'h0000;
            14'h3408: oData <= 16'h0000;
            14'h3409: oData <= 16'h0000;
            14'h340a: oData <= 16'h0000;
            14'h340b: oData <= 16'h0000;
            14'h340c: oData <= 16'h0000;
            14'h340d: oData <= 16'h0000;
            14'h340e: oData <= 16'h0000;
            14'h340f: oData <= 16'h0000;
            14'h3410: oData <= 16'h0000;
            14'h3411: oData <= 16'h0000;
            14'h3412: oData <= 16'h0000;
            14'h3413: oData <= 16'h0000;
            14'h3414: oData <= 16'h0000;
            14'h3415: oData <= 16'h0000;
            14'h3416: oData <= 16'h0000;
            14'h3417: oData <= 16'h0000;
            14'h3418: oData <= 16'h0000;
            14'h3419: oData <= 16'h0000;
            14'h341a: oData <= 16'h0000;
            14'h341b: oData <= 16'h0000;
            14'h341c: oData <= 16'h0000;
            14'h341d: oData <= 16'h0000;
            14'h341e: oData <= 16'h0000;
            14'h341f: oData <= 16'h0000;
            14'h3420: oData <= 16'h0000;
            14'h3421: oData <= 16'h0000;
            14'h3422: oData <= 16'h0000;
            14'h3423: oData <= 16'h0000;
            14'h3424: oData <= 16'h0000;
            14'h3425: oData <= 16'h0000;
            14'h3426: oData <= 16'h0000;
            14'h3427: oData <= 16'h0000;
            14'h3428: oData <= 16'h0000;
            14'h3429: oData <= 16'h0000;
            14'h342a: oData <= 16'h0000;
            14'h342b: oData <= 16'h0000;
            14'h342c: oData <= 16'h0000;
            14'h342d: oData <= 16'h0000;
            14'h342e: oData <= 16'h0000;
            14'h342f: oData <= 16'h0000;
            14'h3430: oData <= 16'h0000;
            14'h3431: oData <= 16'h0000;
            14'h3432: oData <= 16'h0000;
            14'h3433: oData <= 16'h0000;
            14'h3434: oData <= 16'h0000;
            14'h3435: oData <= 16'h0000;
            14'h3436: oData <= 16'h0000;
            14'h3437: oData <= 16'h0000;
            14'h3438: oData <= 16'h0000;
            14'h3439: oData <= 16'h0000;
            14'h343a: oData <= 16'h0000;
            14'h343b: oData <= 16'h0000;
            14'h343c: oData <= 16'h0000;
            14'h343d: oData <= 16'h0000;
            14'h343e: oData <= 16'h0000;
            14'h343f: oData <= 16'h0000;
            14'h3440: oData <= 16'h0000;
            14'h3441: oData <= 16'h0000;
            14'h3442: oData <= 16'h0000;
            14'h3443: oData <= 16'h0000;
            14'h3444: oData <= 16'h0000;
            14'h3445: oData <= 16'h0000;
            14'h3446: oData <= 16'h0000;
            14'h3447: oData <= 16'h0000;
            14'h3448: oData <= 16'h0000;
            14'h3449: oData <= 16'h0000;
            14'h344a: oData <= 16'h0000;
            14'h344b: oData <= 16'h0000;
            14'h344c: oData <= 16'h0000;
            14'h344d: oData <= 16'h0000;
            14'h344e: oData <= 16'h0000;
            14'h344f: oData <= 16'h0000;
            14'h3450: oData <= 16'h0000;
            14'h3451: oData <= 16'h0000;
            14'h3452: oData <= 16'h0000;
            14'h3453: oData <= 16'h0000;
            14'h3454: oData <= 16'h0000;
            14'h3455: oData <= 16'h0000;
            14'h3456: oData <= 16'h0000;
            14'h3457: oData <= 16'h0000;
            14'h3458: oData <= 16'h0000;
            14'h3459: oData <= 16'h0000;
            14'h345a: oData <= 16'h0000;
            14'h345b: oData <= 16'h0000;
            14'h345c: oData <= 16'h0000;
            14'h345d: oData <= 16'h0000;
            14'h345e: oData <= 16'h0000;
            14'h345f: oData <= 16'h0000;
            14'h3460: oData <= 16'h0000;
            14'h3461: oData <= 16'h0000;
            14'h3462: oData <= 16'h0000;
            14'h3463: oData <= 16'h0000;
            14'h3464: oData <= 16'h0000;
            14'h3465: oData <= 16'h0000;
            14'h3466: oData <= 16'h0000;
            14'h3467: oData <= 16'h0000;
            14'h3468: oData <= 16'h0000;
            14'h3469: oData <= 16'h0000;
            14'h346a: oData <= 16'h0000;
            14'h346b: oData <= 16'h0000;
            14'h346c: oData <= 16'h0000;
            14'h346d: oData <= 16'h0000;
            14'h346e: oData <= 16'h0000;
            14'h346f: oData <= 16'h0000;
            14'h3470: oData <= 16'h0000;
            14'h3471: oData <= 16'h0000;
            14'h3472: oData <= 16'h0000;
            14'h3473: oData <= 16'h0000;
            14'h3474: oData <= 16'h0000;
            14'h3475: oData <= 16'h0000;
            14'h3476: oData <= 16'h0000;
            14'h3477: oData <= 16'h0000;
            14'h3478: oData <= 16'h0000;
            14'h3479: oData <= 16'h0000;
            14'h347a: oData <= 16'h0000;
            14'h347b: oData <= 16'h0000;
            14'h347c: oData <= 16'h0000;
            14'h347d: oData <= 16'h0000;
            14'h347e: oData <= 16'h0000;
            14'h347f: oData <= 16'h0000;
            14'h3480: oData <= 16'h0000;
            14'h3481: oData <= 16'h0000;
            14'h3482: oData <= 16'h0000;
            14'h3483: oData <= 16'h0000;
            14'h3484: oData <= 16'h0000;
            14'h3485: oData <= 16'h0000;
            14'h3486: oData <= 16'h0000;
            14'h3487: oData <= 16'h0000;
            14'h3488: oData <= 16'h0000;
            14'h3489: oData <= 16'h0000;
            14'h348a: oData <= 16'h0000;
            14'h348b: oData <= 16'h0000;
            14'h348c: oData <= 16'h0000;
            14'h348d: oData <= 16'h0000;
            14'h348e: oData <= 16'h0000;
            14'h348f: oData <= 16'h0000;
            14'h3490: oData <= 16'h0000;
            14'h3491: oData <= 16'h0000;
            14'h3492: oData <= 16'h0000;
            14'h3493: oData <= 16'h0000;
            14'h3494: oData <= 16'h0000;
            14'h3495: oData <= 16'h0000;
            14'h3496: oData <= 16'h0000;
            14'h3497: oData <= 16'h0000;
            14'h3498: oData <= 16'h0000;
            14'h3499: oData <= 16'h0000;
            14'h349a: oData <= 16'h0000;
            14'h349b: oData <= 16'h0000;
            14'h349c: oData <= 16'h0000;
            14'h349d: oData <= 16'h0000;
            14'h349e: oData <= 16'h0000;
            14'h349f: oData <= 16'h0000;
            14'h34a0: oData <= 16'h0000;
            14'h34a1: oData <= 16'h0000;
            14'h34a2: oData <= 16'h0000;
            14'h34a3: oData <= 16'h0000;
            14'h34a4: oData <= 16'h0000;
            14'h34a5: oData <= 16'h0000;
            14'h34a6: oData <= 16'h0000;
            14'h34a7: oData <= 16'h0000;
            14'h34a8: oData <= 16'h0000;
            14'h34a9: oData <= 16'h0000;
            14'h34aa: oData <= 16'h0000;
            14'h34ab: oData <= 16'h0000;
            14'h34ac: oData <= 16'h0000;
            14'h34ad: oData <= 16'h0000;
            14'h34ae: oData <= 16'h0000;
            14'h34af: oData <= 16'h0000;
            14'h34b0: oData <= 16'h0000;
            14'h34b1: oData <= 16'h0000;
            14'h34b2: oData <= 16'h0000;
            14'h34b3: oData <= 16'h0000;
            14'h34b4: oData <= 16'h0000;
            14'h34b5: oData <= 16'h0000;
            14'h34b6: oData <= 16'h0000;
            14'h34b7: oData <= 16'h0000;
            14'h34b8: oData <= 16'h0000;
            14'h34b9: oData <= 16'h0000;
            14'h34ba: oData <= 16'h0000;
            14'h34bb: oData <= 16'h0000;
            14'h34bc: oData <= 16'h0000;
            14'h34bd: oData <= 16'h0000;
            14'h34be: oData <= 16'h0000;
            14'h34bf: oData <= 16'h0000;
            14'h34c0: oData <= 16'h0000;
            14'h34c1: oData <= 16'h0000;
            14'h34c2: oData <= 16'h0000;
            14'h34c3: oData <= 16'h0000;
            14'h34c4: oData <= 16'h0000;
            14'h34c5: oData <= 16'h0000;
            14'h34c6: oData <= 16'h0000;
            14'h34c7: oData <= 16'h0000;
            14'h34c8: oData <= 16'h0000;
            14'h34c9: oData <= 16'h0000;
            14'h34ca: oData <= 16'h0000;
            14'h34cb: oData <= 16'h0000;
            14'h34cc: oData <= 16'h0000;
            14'h34cd: oData <= 16'h0000;
            14'h34ce: oData <= 16'h0000;
            14'h34cf: oData <= 16'h0000;
            14'h34d0: oData <= 16'h0000;
            14'h34d1: oData <= 16'h0000;
            14'h34d2: oData <= 16'h0000;
            14'h34d3: oData <= 16'h0000;
            14'h34d4: oData <= 16'h0000;
            14'h34d5: oData <= 16'h0000;
            14'h34d6: oData <= 16'h0000;
            14'h34d7: oData <= 16'h0000;
            14'h34d8: oData <= 16'h0000;
            14'h34d9: oData <= 16'h0000;
            14'h34da: oData <= 16'h0000;
            14'h34db: oData <= 16'h0000;
            14'h34dc: oData <= 16'h0000;
            14'h34dd: oData <= 16'h0000;
            14'h34de: oData <= 16'h0000;
            14'h34df: oData <= 16'h0000;
            14'h34e0: oData <= 16'h0000;
            14'h34e1: oData <= 16'h0000;
            14'h34e2: oData <= 16'h0000;
            14'h34e3: oData <= 16'h0000;
            14'h34e4: oData <= 16'h0000;
            14'h34e5: oData <= 16'h0000;
            14'h34e6: oData <= 16'h0000;
            14'h34e7: oData <= 16'h0000;
            14'h34e8: oData <= 16'h0000;
            14'h34e9: oData <= 16'h0000;
            14'h34ea: oData <= 16'h0000;
            14'h34eb: oData <= 16'h0000;
            14'h34ec: oData <= 16'h0000;
            14'h34ed: oData <= 16'h0000;
            14'h34ee: oData <= 16'h0000;
            14'h34ef: oData <= 16'h0000;
            14'h34f0: oData <= 16'h0000;
            14'h34f1: oData <= 16'h0000;
            14'h34f2: oData <= 16'h0000;
            14'h34f3: oData <= 16'h0000;
            14'h34f4: oData <= 16'h0000;
            14'h34f5: oData <= 16'h0000;
            14'h34f6: oData <= 16'h0000;
            14'h34f7: oData <= 16'h0000;
            14'h34f8: oData <= 16'h0000;
            14'h34f9: oData <= 16'h0000;
            14'h34fa: oData <= 16'h0000;
            14'h34fb: oData <= 16'h0000;
            14'h34fc: oData <= 16'h0000;
            14'h34fd: oData <= 16'h0000;
            14'h34fe: oData <= 16'h0000;
            14'h34ff: oData <= 16'h0000;
            14'h3500: oData <= 16'h0000;
            14'h3501: oData <= 16'h0000;
            14'h3502: oData <= 16'h0000;
            14'h3503: oData <= 16'h0000;
            14'h3504: oData <= 16'h0000;
            14'h3505: oData <= 16'h0000;
            14'h3506: oData <= 16'h0000;
            14'h3507: oData <= 16'h0000;
            14'h3508: oData <= 16'h0000;
            14'h3509: oData <= 16'h0000;
            14'h350a: oData <= 16'h0000;
            14'h350b: oData <= 16'h0000;
            14'h350c: oData <= 16'h0000;
            14'h350d: oData <= 16'h0000;
            14'h350e: oData <= 16'h0000;
            14'h350f: oData <= 16'h0000;
            14'h3510: oData <= 16'h0000;
            14'h3511: oData <= 16'h0000;
            14'h3512: oData <= 16'h0000;
            14'h3513: oData <= 16'h0000;
            14'h3514: oData <= 16'h0000;
            14'h3515: oData <= 16'h0000;
            14'h3516: oData <= 16'h0000;
            14'h3517: oData <= 16'h0000;
            14'h3518: oData <= 16'h0000;
            14'h3519: oData <= 16'h0000;
            14'h351a: oData <= 16'h0000;
            14'h351b: oData <= 16'h0000;
            14'h351c: oData <= 16'h0000;
            14'h351d: oData <= 16'h0000;
            14'h351e: oData <= 16'h0000;
            14'h351f: oData <= 16'h0000;
            14'h3520: oData <= 16'h0000;
            14'h3521: oData <= 16'h0000;
            14'h3522: oData <= 16'h0000;
            14'h3523: oData <= 16'h0000;
            14'h3524: oData <= 16'h0000;
            14'h3525: oData <= 16'h0000;
            14'h3526: oData <= 16'h0000;
            14'h3527: oData <= 16'h0000;
            14'h3528: oData <= 16'h0000;
            14'h3529: oData <= 16'h0000;
            14'h352a: oData <= 16'h0000;
            14'h352b: oData <= 16'h0000;
            14'h352c: oData <= 16'h0000;
            14'h352d: oData <= 16'h0000;
            14'h352e: oData <= 16'h0000;
            14'h352f: oData <= 16'h0000;
            14'h3530: oData <= 16'h0000;
            14'h3531: oData <= 16'h0000;
            14'h3532: oData <= 16'h0000;
            14'h3533: oData <= 16'h0000;
            14'h3534: oData <= 16'h0000;
            14'h3535: oData <= 16'h0000;
            14'h3536: oData <= 16'h0000;
            14'h3537: oData <= 16'h0000;
            14'h3538: oData <= 16'h0000;
            14'h3539: oData <= 16'h0000;
            14'h353a: oData <= 16'h0000;
            14'h353b: oData <= 16'h0000;
            14'h353c: oData <= 16'h0000;
            14'h353d: oData <= 16'h0000;
            14'h353e: oData <= 16'h0000;
            14'h353f: oData <= 16'h0000;
            14'h3540: oData <= 16'h0000;
            14'h3541: oData <= 16'h0000;
            14'h3542: oData <= 16'h0000;
            14'h3543: oData <= 16'h0000;
            14'h3544: oData <= 16'h0000;
            14'h3545: oData <= 16'h0000;
            14'h3546: oData <= 16'h0000;
            14'h3547: oData <= 16'h0000;
            14'h3548: oData <= 16'h0000;
            14'h3549: oData <= 16'h0000;
            14'h354a: oData <= 16'h0000;
            14'h354b: oData <= 16'h0000;
            14'h354c: oData <= 16'h0000;
            14'h354d: oData <= 16'h0000;
            14'h354e: oData <= 16'h0000;
            14'h354f: oData <= 16'h0000;
            14'h3550: oData <= 16'h0000;
            14'h3551: oData <= 16'h0000;
            14'h3552: oData <= 16'h0000;
            14'h3553: oData <= 16'h0000;
            14'h3554: oData <= 16'h0000;
            14'h3555: oData <= 16'h0000;
            14'h3556: oData <= 16'h0000;
            14'h3557: oData <= 16'h0000;
            14'h3558: oData <= 16'h0000;
            14'h3559: oData <= 16'h0000;
            14'h355a: oData <= 16'h0000;
            14'h355b: oData <= 16'h0000;
            14'h355c: oData <= 16'h0000;
            14'h355d: oData <= 16'h0000;
            14'h355e: oData <= 16'h0000;
            14'h355f: oData <= 16'h0000;
            14'h3560: oData <= 16'h0000;
            14'h3561: oData <= 16'h0000;
            14'h3562: oData <= 16'h0000;
            14'h3563: oData <= 16'h0000;
            14'h3564: oData <= 16'h0000;
            14'h3565: oData <= 16'h0000;
            14'h3566: oData <= 16'h0000;
            14'h3567: oData <= 16'h0000;
            14'h3568: oData <= 16'h0000;
            14'h3569: oData <= 16'h0000;
            14'h356a: oData <= 16'h0000;
            14'h356b: oData <= 16'h0000;
            14'h356c: oData <= 16'h0000;
            14'h356d: oData <= 16'h0000;
            14'h356e: oData <= 16'h0000;
            14'h356f: oData <= 16'h0000;
            14'h3570: oData <= 16'h0000;
            14'h3571: oData <= 16'h0000;
            14'h3572: oData <= 16'h0000;
            14'h3573: oData <= 16'h0000;
            14'h3574: oData <= 16'h0000;
            14'h3575: oData <= 16'h0000;
            14'h3576: oData <= 16'h0000;
            14'h3577: oData <= 16'h0000;
            14'h3578: oData <= 16'h0000;
            14'h3579: oData <= 16'h0000;
            14'h357a: oData <= 16'h0000;
            14'h357b: oData <= 16'h0000;
            14'h357c: oData <= 16'h0000;
            14'h357d: oData <= 16'h0000;
            14'h357e: oData <= 16'h0000;
            14'h357f: oData <= 16'h0000;
            14'h3580: oData <= 16'h0000;
            14'h3581: oData <= 16'h0000;
            14'h3582: oData <= 16'h0000;
            14'h3583: oData <= 16'h0000;
            14'h3584: oData <= 16'h0000;
            14'h3585: oData <= 16'h0000;
            14'h3586: oData <= 16'h0000;
            14'h3587: oData <= 16'h0000;
            14'h3588: oData <= 16'h0000;
            14'h3589: oData <= 16'h0000;
            14'h358a: oData <= 16'h0000;
            14'h358b: oData <= 16'h0000;
            14'h358c: oData <= 16'h0000;
            14'h358d: oData <= 16'h0000;
            14'h358e: oData <= 16'h0000;
            14'h358f: oData <= 16'h0000;
            14'h3590: oData <= 16'h0000;
            14'h3591: oData <= 16'h0000;
            14'h3592: oData <= 16'h0000;
            14'h3593: oData <= 16'h0000;
            14'h3594: oData <= 16'h0000;
            14'h3595: oData <= 16'h0000;
            14'h3596: oData <= 16'h0000;
            14'h3597: oData <= 16'h0000;
            14'h3598: oData <= 16'h0000;
            14'h3599: oData <= 16'h0000;
            14'h359a: oData <= 16'h0000;
            14'h359b: oData <= 16'h0000;
            14'h359c: oData <= 16'h0000;
            14'h359d: oData <= 16'h0000;
            14'h359e: oData <= 16'h0000;
            14'h359f: oData <= 16'h0000;
            14'h35a0: oData <= 16'h0000;
            14'h35a1: oData <= 16'h0000;
            14'h35a2: oData <= 16'h0000;
            14'h35a3: oData <= 16'h0000;
            14'h35a4: oData <= 16'h0000;
            14'h35a5: oData <= 16'h0000;
            14'h35a6: oData <= 16'h0000;
            14'h35a7: oData <= 16'h0000;
            14'h35a8: oData <= 16'h0000;
            14'h35a9: oData <= 16'h0000;
            14'h35aa: oData <= 16'h0000;
            14'h35ab: oData <= 16'h0000;
            14'h35ac: oData <= 16'h0000;
            14'h35ad: oData <= 16'h0000;
            14'h35ae: oData <= 16'h0000;
            14'h35af: oData <= 16'h0000;
            14'h35b0: oData <= 16'h0000;
            14'h35b1: oData <= 16'h0000;
            14'h35b2: oData <= 16'h0000;
            14'h35b3: oData <= 16'h0000;
            14'h35b4: oData <= 16'h0000;
            14'h35b5: oData <= 16'h0000;
            14'h35b6: oData <= 16'h0000;
            14'h35b7: oData <= 16'h0000;
            14'h35b8: oData <= 16'h0000;
            14'h35b9: oData <= 16'h0000;
            14'h35ba: oData <= 16'h0000;
            14'h35bb: oData <= 16'h0000;
            14'h35bc: oData <= 16'h0000;
            14'h35bd: oData <= 16'h0000;
            14'h35be: oData <= 16'h0000;
            14'h35bf: oData <= 16'h0000;
            14'h35c0: oData <= 16'h0000;
            14'h35c1: oData <= 16'h0000;
            14'h35c2: oData <= 16'h0000;
            14'h35c3: oData <= 16'h0000;
            14'h35c4: oData <= 16'h0000;
            14'h35c5: oData <= 16'h0000;
            14'h35c6: oData <= 16'h0000;
            14'h35c7: oData <= 16'h0000;
            14'h35c8: oData <= 16'h0000;
            14'h35c9: oData <= 16'h0000;
            14'h35ca: oData <= 16'h0000;
            14'h35cb: oData <= 16'h0000;
            14'h35cc: oData <= 16'h0000;
            14'h35cd: oData <= 16'h0000;
            14'h35ce: oData <= 16'h0000;
            14'h35cf: oData <= 16'h0000;
            14'h35d0: oData <= 16'h0000;
            14'h35d1: oData <= 16'h0000;
            14'h35d2: oData <= 16'h0000;
            14'h35d3: oData <= 16'h0000;
            14'h35d4: oData <= 16'h0000;
            14'h35d5: oData <= 16'h0000;
            14'h35d6: oData <= 16'h0000;
            14'h35d7: oData <= 16'h0000;
            14'h35d8: oData <= 16'h0000;
            14'h35d9: oData <= 16'h0000;
            14'h35da: oData <= 16'h0000;
            14'h35db: oData <= 16'h0000;
            14'h35dc: oData <= 16'h0000;
            14'h35dd: oData <= 16'h0000;
            14'h35de: oData <= 16'h0000;
            14'h35df: oData <= 16'h0000;
            14'h35e0: oData <= 16'h0000;
            14'h35e1: oData <= 16'h0000;
            14'h35e2: oData <= 16'h0000;
            14'h35e3: oData <= 16'h0000;
            14'h35e4: oData <= 16'h0000;
            14'h35e5: oData <= 16'h0000;
            14'h35e6: oData <= 16'h0000;
            14'h35e7: oData <= 16'h0000;
            14'h35e8: oData <= 16'h0000;
            14'h35e9: oData <= 16'h0000;
            14'h35ea: oData <= 16'h0000;
            14'h35eb: oData <= 16'h0000;
            14'h35ec: oData <= 16'h0000;
            14'h35ed: oData <= 16'h0000;
            14'h35ee: oData <= 16'h0000;
            14'h35ef: oData <= 16'h0000;
            14'h35f0: oData <= 16'h0000;
            14'h35f1: oData <= 16'h0000;
            14'h35f2: oData <= 16'h0000;
            14'h35f3: oData <= 16'h0000;
            14'h35f4: oData <= 16'h0000;
            14'h35f5: oData <= 16'h0000;
            14'h35f6: oData <= 16'h0000;
            14'h35f7: oData <= 16'h0000;
            14'h35f8: oData <= 16'h0000;
            14'h35f9: oData <= 16'h0000;
            14'h35fa: oData <= 16'h0000;
            14'h35fb: oData <= 16'h0000;
            14'h35fc: oData <= 16'h0000;
            14'h35fd: oData <= 16'h0000;
            14'h35fe: oData <= 16'h0000;
            14'h35ff: oData <= 16'h0000;
            14'h3600: oData <= 16'h0000;
            14'h3601: oData <= 16'h0000;
            14'h3602: oData <= 16'h0000;
            14'h3603: oData <= 16'h0000;
            14'h3604: oData <= 16'h0000;
            14'h3605: oData <= 16'h0000;
            14'h3606: oData <= 16'h0000;
            14'h3607: oData <= 16'h0000;
            14'h3608: oData <= 16'h0000;
            14'h3609: oData <= 16'h0000;
            14'h360a: oData <= 16'h0000;
            14'h360b: oData <= 16'h0000;
            14'h360c: oData <= 16'h0000;
            14'h360d: oData <= 16'h0000;
            14'h360e: oData <= 16'h0000;
            14'h360f: oData <= 16'h0000;
            14'h3610: oData <= 16'h0000;
            14'h3611: oData <= 16'h0000;
            14'h3612: oData <= 16'h0000;
            14'h3613: oData <= 16'h0000;
            14'h3614: oData <= 16'h0000;
            14'h3615: oData <= 16'h0000;
            14'h3616: oData <= 16'h0000;
            14'h3617: oData <= 16'h0000;
            14'h3618: oData <= 16'h0000;
            14'h3619: oData <= 16'h0000;
            14'h361a: oData <= 16'h0000;
            14'h361b: oData <= 16'h0000;
            14'h361c: oData <= 16'h0000;
            14'h361d: oData <= 16'h0000;
            14'h361e: oData <= 16'h0000;
            14'h361f: oData <= 16'h0000;
            14'h3620: oData <= 16'h0000;
            14'h3621: oData <= 16'h0000;
            14'h3622: oData <= 16'h0000;
            14'h3623: oData <= 16'h0000;
            14'h3624: oData <= 16'h0000;
            14'h3625: oData <= 16'h0000;
            14'h3626: oData <= 16'h0000;
            14'h3627: oData <= 16'h0000;
            14'h3628: oData <= 16'h0000;
            14'h3629: oData <= 16'h0000;
            14'h362a: oData <= 16'h0000;
            14'h362b: oData <= 16'h0000;
            14'h362c: oData <= 16'h0000;
            14'h362d: oData <= 16'h0000;
            14'h362e: oData <= 16'h0000;
            14'h362f: oData <= 16'h0000;
            14'h3630: oData <= 16'h0000;
            14'h3631: oData <= 16'h0000;
            14'h3632: oData <= 16'h0000;
            14'h3633: oData <= 16'h0000;
            14'h3634: oData <= 16'h0000;
            14'h3635: oData <= 16'h0000;
            14'h3636: oData <= 16'h0000;
            14'h3637: oData <= 16'h0000;
            14'h3638: oData <= 16'h0000;
            14'h3639: oData <= 16'h0000;
            14'h363a: oData <= 16'h0000;
            14'h363b: oData <= 16'h0000;
            14'h363c: oData <= 16'h0000;
            14'h363d: oData <= 16'h0000;
            14'h363e: oData <= 16'h0000;
            14'h363f: oData <= 16'h0000;
            14'h3640: oData <= 16'h0000;
            14'h3641: oData <= 16'h0000;
            14'h3642: oData <= 16'h0000;
            14'h3643: oData <= 16'h0000;
            14'h3644: oData <= 16'h0000;
            14'h3645: oData <= 16'h0000;
            14'h3646: oData <= 16'h0000;
            14'h3647: oData <= 16'h0000;
            14'h3648: oData <= 16'h0000;
            14'h3649: oData <= 16'h0000;
            14'h364a: oData <= 16'h0000;
            14'h364b: oData <= 16'h0000;
            14'h364c: oData <= 16'h0000;
            14'h364d: oData <= 16'h0000;
            14'h364e: oData <= 16'h0000;
            14'h364f: oData <= 16'h0000;
            14'h3650: oData <= 16'h0000;
            14'h3651: oData <= 16'h0000;
            14'h3652: oData <= 16'h0000;
            14'h3653: oData <= 16'h0000;
            14'h3654: oData <= 16'h0000;
            14'h3655: oData <= 16'h0000;
            14'h3656: oData <= 16'h0000;
            14'h3657: oData <= 16'h0000;
            14'h3658: oData <= 16'h0000;
            14'h3659: oData <= 16'h0000;
            14'h365a: oData <= 16'h0000;
            14'h365b: oData <= 16'h0000;
            14'h365c: oData <= 16'h0000;
            14'h365d: oData <= 16'h0000;
            14'h365e: oData <= 16'h0000;
            14'h365f: oData <= 16'h0000;
            14'h3660: oData <= 16'h0000;
            14'h3661: oData <= 16'h0000;
            14'h3662: oData <= 16'h0000;
            14'h3663: oData <= 16'h0000;
            14'h3664: oData <= 16'h0000;
            14'h3665: oData <= 16'h0000;
            14'h3666: oData <= 16'h0000;
            14'h3667: oData <= 16'h0000;
            14'h3668: oData <= 16'h0000;
            14'h3669: oData <= 16'h0000;
            14'h366a: oData <= 16'h0000;
            14'h366b: oData <= 16'h0000;
            14'h366c: oData <= 16'h0000;
            14'h366d: oData <= 16'h0000;
            14'h366e: oData <= 16'h0000;
            14'h366f: oData <= 16'h0000;
            14'h3670: oData <= 16'h0000;
            14'h3671: oData <= 16'h0000;
            14'h3672: oData <= 16'h0000;
            14'h3673: oData <= 16'h0000;
            14'h3674: oData <= 16'h0000;
            14'h3675: oData <= 16'h0000;
            14'h3676: oData <= 16'h0000;
            14'h3677: oData <= 16'h0000;
            14'h3678: oData <= 16'h0000;
            14'h3679: oData <= 16'h0000;
            14'h367a: oData <= 16'h0000;
            14'h367b: oData <= 16'h0000;
            14'h367c: oData <= 16'h0000;
            14'h367d: oData <= 16'h0000;
            14'h367e: oData <= 16'h0000;
            14'h367f: oData <= 16'h0000;
            14'h3680: oData <= 16'h0000;
            14'h3681: oData <= 16'h0000;
            14'h3682: oData <= 16'h0000;
            14'h3683: oData <= 16'h0000;
            14'h3684: oData <= 16'h0000;
            14'h3685: oData <= 16'h0000;
            14'h3686: oData <= 16'h0000;
            14'h3687: oData <= 16'h0000;
            14'h3688: oData <= 16'h0000;
            14'h3689: oData <= 16'h0000;
            14'h368a: oData <= 16'h0000;
            14'h368b: oData <= 16'h0000;
            14'h368c: oData <= 16'h0000;
            14'h368d: oData <= 16'h0000;
            14'h368e: oData <= 16'h0000;
            14'h368f: oData <= 16'h0000;
            14'h3690: oData <= 16'h0000;
            14'h3691: oData <= 16'h0000;
            14'h3692: oData <= 16'h0000;
            14'h3693: oData <= 16'h0000;
            14'h3694: oData <= 16'h0000;
            14'h3695: oData <= 16'h0000;
            14'h3696: oData <= 16'h0000;
            14'h3697: oData <= 16'h0000;
            14'h3698: oData <= 16'h0000;
            14'h3699: oData <= 16'h0000;
            14'h369a: oData <= 16'h0000;
            14'h369b: oData <= 16'h0000;
            14'h369c: oData <= 16'h0000;
            14'h369d: oData <= 16'h0000;
            14'h369e: oData <= 16'h0000;
            14'h369f: oData <= 16'h0000;
            14'h36a0: oData <= 16'h0000;
            14'h36a1: oData <= 16'h0000;
            14'h36a2: oData <= 16'h0000;
            14'h36a3: oData <= 16'h0000;
            14'h36a4: oData <= 16'h0000;
            14'h36a5: oData <= 16'h0000;
            14'h36a6: oData <= 16'h0000;
            14'h36a7: oData <= 16'h0000;
            14'h36a8: oData <= 16'h0000;
            14'h36a9: oData <= 16'h0000;
            14'h36aa: oData <= 16'h0000;
            14'h36ab: oData <= 16'h0000;
            14'h36ac: oData <= 16'h0000;
            14'h36ad: oData <= 16'h0000;
            14'h36ae: oData <= 16'h0000;
            14'h36af: oData <= 16'h0000;
            14'h36b0: oData <= 16'h0000;
            14'h36b1: oData <= 16'h0000;
            14'h36b2: oData <= 16'h0000;
            14'h36b3: oData <= 16'h0000;
            14'h36b4: oData <= 16'h0000;
            14'h36b5: oData <= 16'h0000;
            14'h36b6: oData <= 16'h0000;
            14'h36b7: oData <= 16'h0000;
            14'h36b8: oData <= 16'h0000;
            14'h36b9: oData <= 16'h0000;
            14'h36ba: oData <= 16'h0000;
            14'h36bb: oData <= 16'h0000;
            14'h36bc: oData <= 16'h0000;
            14'h36bd: oData <= 16'h0000;
            14'h36be: oData <= 16'h0000;
            14'h36bf: oData <= 16'h0000;
            14'h36c0: oData <= 16'h0000;
            14'h36c1: oData <= 16'h0000;
            14'h36c2: oData <= 16'h0000;
            14'h36c3: oData <= 16'h0000;
            14'h36c4: oData <= 16'h0000;
            14'h36c5: oData <= 16'h0000;
            14'h36c6: oData <= 16'h0000;
            14'h36c7: oData <= 16'h0000;
            14'h36c8: oData <= 16'h0000;
            14'h36c9: oData <= 16'h0000;
            14'h36ca: oData <= 16'h0000;
            14'h36cb: oData <= 16'h0000;
            14'h36cc: oData <= 16'h0000;
            14'h36cd: oData <= 16'h0000;
            14'h36ce: oData <= 16'h0000;
            14'h36cf: oData <= 16'h0000;
            14'h36d0: oData <= 16'h0000;
            14'h36d1: oData <= 16'h0000;
            14'h36d2: oData <= 16'h0000;
            14'h36d3: oData <= 16'h0000;
            14'h36d4: oData <= 16'h0000;
            14'h36d5: oData <= 16'h0000;
            14'h36d6: oData <= 16'h0000;
            14'h36d7: oData <= 16'h0000;
            14'h36d8: oData <= 16'h0000;
            14'h36d9: oData <= 16'h0000;
            14'h36da: oData <= 16'h0000;
            14'h36db: oData <= 16'h0000;
            14'h36dc: oData <= 16'h0000;
            14'h36dd: oData <= 16'h0000;
            14'h36de: oData <= 16'h0000;
            14'h36df: oData <= 16'h0000;
            14'h36e0: oData <= 16'h0000;
            14'h36e1: oData <= 16'h0000;
            14'h36e2: oData <= 16'h0000;
            14'h36e3: oData <= 16'h0000;
            14'h36e4: oData <= 16'h0000;
            14'h36e5: oData <= 16'h0000;
            14'h36e6: oData <= 16'h0000;
            14'h36e7: oData <= 16'h0000;
            14'h36e8: oData <= 16'h0000;
            14'h36e9: oData <= 16'h0000;
            14'h36ea: oData <= 16'h0000;
            14'h36eb: oData <= 16'h0000;
            14'h36ec: oData <= 16'h0000;
            14'h36ed: oData <= 16'h0000;
            14'h36ee: oData <= 16'h0000;
            14'h36ef: oData <= 16'h0000;
            14'h36f0: oData <= 16'h0000;
            14'h36f1: oData <= 16'h0000;
            14'h36f2: oData <= 16'h0000;
            14'h36f3: oData <= 16'h0000;
            14'h36f4: oData <= 16'h0000;
            14'h36f5: oData <= 16'h0000;
            14'h36f6: oData <= 16'h0000;
            14'h36f7: oData <= 16'h0000;
            14'h36f8: oData <= 16'h0000;
            14'h36f9: oData <= 16'h0000;
            14'h36fa: oData <= 16'h0000;
            14'h36fb: oData <= 16'h0000;
            14'h36fc: oData <= 16'h0000;
            14'h36fd: oData <= 16'h0000;
            14'h36fe: oData <= 16'h0000;
            14'h36ff: oData <= 16'h0000;
            14'h3700: oData <= 16'h0000;
            14'h3701: oData <= 16'h0000;
            14'h3702: oData <= 16'h0000;
            14'h3703: oData <= 16'h0000;
            14'h3704: oData <= 16'h0000;
            14'h3705: oData <= 16'h0000;
            14'h3706: oData <= 16'h0000;
            14'h3707: oData <= 16'h0000;
            14'h3708: oData <= 16'h0000;
            14'h3709: oData <= 16'h0000;
            14'h370a: oData <= 16'h0000;
            14'h370b: oData <= 16'h0000;
            14'h370c: oData <= 16'h0000;
            14'h370d: oData <= 16'h0000;
            14'h370e: oData <= 16'h0000;
            14'h370f: oData <= 16'h0000;
            14'h3710: oData <= 16'h0000;
            14'h3711: oData <= 16'h0000;
            14'h3712: oData <= 16'h0000;
            14'h3713: oData <= 16'h0000;
            14'h3714: oData <= 16'h0000;
            14'h3715: oData <= 16'h0000;
            14'h3716: oData <= 16'h0000;
            14'h3717: oData <= 16'h0000;
            14'h3718: oData <= 16'h0000;
            14'h3719: oData <= 16'h0000;
            14'h371a: oData <= 16'h0000;
            14'h371b: oData <= 16'h0000;
            14'h371c: oData <= 16'h0000;
            14'h371d: oData <= 16'h0000;
            14'h371e: oData <= 16'h0000;
            14'h371f: oData <= 16'h0000;
            14'h3720: oData <= 16'h0000;
            14'h3721: oData <= 16'h0000;
            14'h3722: oData <= 16'h0000;
            14'h3723: oData <= 16'h0000;
            14'h3724: oData <= 16'h0000;
            14'h3725: oData <= 16'h0000;
            14'h3726: oData <= 16'h0000;
            14'h3727: oData <= 16'h0000;
            14'h3728: oData <= 16'h0000;
            14'h3729: oData <= 16'h0000;
            14'h372a: oData <= 16'h0000;
            14'h372b: oData <= 16'h0000;
            14'h372c: oData <= 16'h0000;
            14'h372d: oData <= 16'h0000;
            14'h372e: oData <= 16'h0000;
            14'h372f: oData <= 16'h0000;
            14'h3730: oData <= 16'h0000;
            14'h3731: oData <= 16'h0000;
            14'h3732: oData <= 16'h0000;
            14'h3733: oData <= 16'h0000;
            14'h3734: oData <= 16'h0000;
            14'h3735: oData <= 16'h0000;
            14'h3736: oData <= 16'h0000;
            14'h3737: oData <= 16'h0000;
            14'h3738: oData <= 16'h0000;
            14'h3739: oData <= 16'h0000;
            14'h373a: oData <= 16'h0000;
            14'h373b: oData <= 16'h0000;
            14'h373c: oData <= 16'h0000;
            14'h373d: oData <= 16'h0000;
            14'h373e: oData <= 16'h0000;
            14'h373f: oData <= 16'h0000;
            14'h3740: oData <= 16'h0000;
            14'h3741: oData <= 16'h0000;
            14'h3742: oData <= 16'h0000;
            14'h3743: oData <= 16'h0000;
            14'h3744: oData <= 16'h0000;
            14'h3745: oData <= 16'h0000;
            14'h3746: oData <= 16'h0000;
            14'h3747: oData <= 16'h0000;
            14'h3748: oData <= 16'h0000;
            14'h3749: oData <= 16'h0000;
            14'h374a: oData <= 16'h0000;
            14'h374b: oData <= 16'h0000;
            14'h374c: oData <= 16'h0000;
            14'h374d: oData <= 16'h0000;
            14'h374e: oData <= 16'h0000;
            14'h374f: oData <= 16'h0000;
            14'h3750: oData <= 16'h0000;
            14'h3751: oData <= 16'h0000;
            14'h3752: oData <= 16'h0000;
            14'h3753: oData <= 16'h0000;
            14'h3754: oData <= 16'h0000;
            14'h3755: oData <= 16'h0000;
            14'h3756: oData <= 16'h0000;
            14'h3757: oData <= 16'h0000;
            14'h3758: oData <= 16'h0000;
            14'h3759: oData <= 16'h0000;
            14'h375a: oData <= 16'h0000;
            14'h375b: oData <= 16'h0000;
            14'h375c: oData <= 16'h0000;
            14'h375d: oData <= 16'h0000;
            14'h375e: oData <= 16'h0000;
            14'h375f: oData <= 16'h0000;
            14'h3760: oData <= 16'h0000;
            14'h3761: oData <= 16'h0000;
            14'h3762: oData <= 16'h0000;
            14'h3763: oData <= 16'h0000;
            14'h3764: oData <= 16'h0000;
            14'h3765: oData <= 16'h0000;
            14'h3766: oData <= 16'h0000;
            14'h3767: oData <= 16'h0000;
            14'h3768: oData <= 16'h0000;
            14'h3769: oData <= 16'h0000;
            14'h376a: oData <= 16'h0000;
            14'h376b: oData <= 16'h0000;
            14'h376c: oData <= 16'h0000;
            14'h376d: oData <= 16'h0000;
            14'h376e: oData <= 16'h0000;
            14'h376f: oData <= 16'h0000;
            14'h3770: oData <= 16'h0000;
            14'h3771: oData <= 16'h0000;
            14'h3772: oData <= 16'h0000;
            14'h3773: oData <= 16'h0000;
            14'h3774: oData <= 16'h0000;
            14'h3775: oData <= 16'h0000;
            14'h3776: oData <= 16'h0000;
            14'h3777: oData <= 16'h0000;
            14'h3778: oData <= 16'h0000;
            14'h3779: oData <= 16'h0000;
            14'h377a: oData <= 16'h0000;
            14'h377b: oData <= 16'h0000;
            14'h377c: oData <= 16'h0000;
            14'h377d: oData <= 16'h0000;
            14'h377e: oData <= 16'h0000;
            14'h377f: oData <= 16'h0000;
            14'h3780: oData <= 16'h0000;
            14'h3781: oData <= 16'h0000;
            14'h3782: oData <= 16'h0000;
            14'h3783: oData <= 16'h0000;
            14'h3784: oData <= 16'h0000;
            14'h3785: oData <= 16'h0000;
            14'h3786: oData <= 16'h0000;
            14'h3787: oData <= 16'h0000;
            14'h3788: oData <= 16'h0000;
            14'h3789: oData <= 16'h0000;
            14'h378a: oData <= 16'h0000;
            14'h378b: oData <= 16'h0000;
            14'h378c: oData <= 16'h0000;
            14'h378d: oData <= 16'h0000;
            14'h378e: oData <= 16'h0000;
            14'h378f: oData <= 16'h0000;
            14'h3790: oData <= 16'h0000;
            14'h3791: oData <= 16'h0000;
            14'h3792: oData <= 16'h0000;
            14'h3793: oData <= 16'h0000;
            14'h3794: oData <= 16'h0000;
            14'h3795: oData <= 16'h0000;
            14'h3796: oData <= 16'h0000;
            14'h3797: oData <= 16'h0000;
            14'h3798: oData <= 16'h0000;
            14'h3799: oData <= 16'h0000;
            14'h379a: oData <= 16'h0000;
            14'h379b: oData <= 16'h0000;
            14'h379c: oData <= 16'h0000;
            14'h379d: oData <= 16'h0000;
            14'h379e: oData <= 16'h0000;
            14'h379f: oData <= 16'h0000;
            14'h37a0: oData <= 16'h0000;
            14'h37a1: oData <= 16'h0000;
            14'h37a2: oData <= 16'h0000;
            14'h37a3: oData <= 16'h0000;
            14'h37a4: oData <= 16'h0000;
            14'h37a5: oData <= 16'h0000;
            14'h37a6: oData <= 16'h0000;
            14'h37a7: oData <= 16'h0000;
            14'h37a8: oData <= 16'h0000;
            14'h37a9: oData <= 16'h0000;
            14'h37aa: oData <= 16'h0000;
            14'h37ab: oData <= 16'h0000;
            14'h37ac: oData <= 16'h0000;
            14'h37ad: oData <= 16'h0000;
            14'h37ae: oData <= 16'h0000;
            14'h37af: oData <= 16'h0000;
            14'h37b0: oData <= 16'h0000;
            14'h37b1: oData <= 16'h0000;
            14'h37b2: oData <= 16'h0000;
            14'h37b3: oData <= 16'h0000;
            14'h37b4: oData <= 16'h0000;
            14'h37b5: oData <= 16'h0000;
            14'h37b6: oData <= 16'h0000;
            14'h37b7: oData <= 16'h0000;
            14'h37b8: oData <= 16'h0000;
            14'h37b9: oData <= 16'h0000;
            14'h37ba: oData <= 16'h0000;
            14'h37bb: oData <= 16'h0000;
            14'h37bc: oData <= 16'h0000;
            14'h37bd: oData <= 16'h0000;
            14'h37be: oData <= 16'h0000;
            14'h37bf: oData <= 16'h0000;
            14'h37c0: oData <= 16'h0000;
            14'h37c1: oData <= 16'h0000;
            14'h37c2: oData <= 16'h0000;
            14'h37c3: oData <= 16'h0000;
            14'h37c4: oData <= 16'h0000;
            14'h37c5: oData <= 16'h0000;
            14'h37c6: oData <= 16'h0000;
            14'h37c7: oData <= 16'h0000;
            14'h37c8: oData <= 16'h0000;
            14'h37c9: oData <= 16'h0000;
            14'h37ca: oData <= 16'h0000;
            14'h37cb: oData <= 16'h0000;
            14'h37cc: oData <= 16'h0000;
            14'h37cd: oData <= 16'h0000;
            14'h37ce: oData <= 16'h0000;
            14'h37cf: oData <= 16'h0000;
            14'h37d0: oData <= 16'h0000;
            14'h37d1: oData <= 16'h0000;
            14'h37d2: oData <= 16'h0000;
            14'h37d3: oData <= 16'h0000;
            14'h37d4: oData <= 16'h0000;
            14'h37d5: oData <= 16'h0000;
            14'h37d6: oData <= 16'h0000;
            14'h37d7: oData <= 16'h0000;
            14'h37d8: oData <= 16'h0000;
            14'h37d9: oData <= 16'h0000;
            14'h37da: oData <= 16'h0000;
            14'h37db: oData <= 16'h0000;
            14'h37dc: oData <= 16'h0000;
            14'h37dd: oData <= 16'h0000;
            14'h37de: oData <= 16'h0000;
            14'h37df: oData <= 16'h0000;
            14'h37e0: oData <= 16'h0000;
            14'h37e1: oData <= 16'h0000;
            14'h37e2: oData <= 16'h0000;
            14'h37e3: oData <= 16'h0000;
            14'h37e4: oData <= 16'h0000;
            14'h37e5: oData <= 16'h0000;
            14'h37e6: oData <= 16'h0000;
            14'h37e7: oData <= 16'h0000;
            14'h37e8: oData <= 16'h0000;
            14'h37e9: oData <= 16'h0000;
            14'h37ea: oData <= 16'h0000;
            14'h37eb: oData <= 16'h0000;
            14'h37ec: oData <= 16'h0000;
            14'h37ed: oData <= 16'h0000;
            14'h37ee: oData <= 16'h0000;
            14'h37ef: oData <= 16'h0000;
            14'h37f0: oData <= 16'h0000;
            14'h37f1: oData <= 16'h0000;
            14'h37f2: oData <= 16'h0000;
            14'h37f3: oData <= 16'h0000;
            14'h37f4: oData <= 16'h0000;
            14'h37f5: oData <= 16'h0000;
            14'h37f6: oData <= 16'h0000;
            14'h37f7: oData <= 16'h0000;
            14'h37f8: oData <= 16'h0000;
            14'h37f9: oData <= 16'h0000;
            14'h37fa: oData <= 16'h0000;
            14'h37fb: oData <= 16'h0000;
            14'h37fc: oData <= 16'h0000;
            14'h37fd: oData <= 16'h0000;
            14'h37fe: oData <= 16'h0000;
            14'h37ff: oData <= 16'h0000;
            14'h3800: oData <= 16'h0000;
            14'h3801: oData <= 16'h0000;
            14'h3802: oData <= 16'h0000;
            14'h3803: oData <= 16'h0000;
            14'h3804: oData <= 16'h0000;
            14'h3805: oData <= 16'h0000;
            14'h3806: oData <= 16'h0000;
            14'h3807: oData <= 16'h0000;
            14'h3808: oData <= 16'h0000;
            14'h3809: oData <= 16'h0000;
            14'h380a: oData <= 16'h0000;
            14'h380b: oData <= 16'h0000;
            14'h380c: oData <= 16'h0000;
            14'h380d: oData <= 16'h0000;
            14'h380e: oData <= 16'h0000;
            14'h380f: oData <= 16'h0000;
            14'h3810: oData <= 16'h0000;
            14'h3811: oData <= 16'h0000;
            14'h3812: oData <= 16'h0000;
            14'h3813: oData <= 16'h0000;
            14'h3814: oData <= 16'h0000;
            14'h3815: oData <= 16'h0000;
            14'h3816: oData <= 16'h0000;
            14'h3817: oData <= 16'h0000;
            14'h3818: oData <= 16'h0000;
            14'h3819: oData <= 16'h0000;
            14'h381a: oData <= 16'h0000;
            14'h381b: oData <= 16'h0000;
            14'h381c: oData <= 16'h0000;
            14'h381d: oData <= 16'h0000;
            14'h381e: oData <= 16'h0000;
            14'h381f: oData <= 16'h0000;
            14'h3820: oData <= 16'h0000;
            14'h3821: oData <= 16'h0000;
            14'h3822: oData <= 16'h0000;
            14'h3823: oData <= 16'h0000;
            14'h3824: oData <= 16'h0000;
            14'h3825: oData <= 16'h0000;
            14'h3826: oData <= 16'h0000;
            14'h3827: oData <= 16'h0000;
            14'h3828: oData <= 16'h0000;
            14'h3829: oData <= 16'h0000;
            14'h382a: oData <= 16'h0000;
            14'h382b: oData <= 16'h0000;
            14'h382c: oData <= 16'h0000;
            14'h382d: oData <= 16'h0000;
            14'h382e: oData <= 16'h0000;
            14'h382f: oData <= 16'h0000;
            14'h3830: oData <= 16'h0000;
            14'h3831: oData <= 16'h0000;
            14'h3832: oData <= 16'h0000;
            14'h3833: oData <= 16'h0000;
            14'h3834: oData <= 16'h0000;
            14'h3835: oData <= 16'h0000;
            14'h3836: oData <= 16'h0000;
            14'h3837: oData <= 16'h0000;
            14'h3838: oData <= 16'h0000;
            14'h3839: oData <= 16'h0000;
            14'h383a: oData <= 16'h0000;
            14'h383b: oData <= 16'h0000;
            14'h383c: oData <= 16'h0000;
            14'h383d: oData <= 16'h0000;
            14'h383e: oData <= 16'h0000;
            14'h383f: oData <= 16'h0000;
            14'h3840: oData <= 16'h0000;
            14'h3841: oData <= 16'h0000;
            14'h3842: oData <= 16'h0000;
            14'h3843: oData <= 16'h0000;
            14'h3844: oData <= 16'h0000;
            14'h3845: oData <= 16'h0000;
            14'h3846: oData <= 16'h0000;
            14'h3847: oData <= 16'h0000;
            14'h3848: oData <= 16'h0000;
            14'h3849: oData <= 16'h0000;
            14'h384a: oData <= 16'h0000;
            14'h384b: oData <= 16'h0000;
            14'h384c: oData <= 16'h0000;
            14'h384d: oData <= 16'h0000;
            14'h384e: oData <= 16'h0000;
            14'h384f: oData <= 16'h0000;
            14'h3850: oData <= 16'h0000;
            14'h3851: oData <= 16'h0000;
            14'h3852: oData <= 16'h0000;
            14'h3853: oData <= 16'h0000;
            14'h3854: oData <= 16'h0000;
            14'h3855: oData <= 16'h0000;
            14'h3856: oData <= 16'h0000;
            14'h3857: oData <= 16'h0000;
            14'h3858: oData <= 16'h0000;
            14'h3859: oData <= 16'h0000;
            14'h385a: oData <= 16'h0000;
            14'h385b: oData <= 16'h0000;
            14'h385c: oData <= 16'h0000;
            14'h385d: oData <= 16'h0000;
            14'h385e: oData <= 16'h0000;
            14'h385f: oData <= 16'h0000;
            14'h3860: oData <= 16'h0000;
            14'h3861: oData <= 16'h0000;
            14'h3862: oData <= 16'h0000;
            14'h3863: oData <= 16'h0000;
            14'h3864: oData <= 16'h0000;
            14'h3865: oData <= 16'h0000;
            14'h3866: oData <= 16'h0000;
            14'h3867: oData <= 16'h0000;
            14'h3868: oData <= 16'h0000;
            14'h3869: oData <= 16'h0000;
            14'h386a: oData <= 16'h0000;
            14'h386b: oData <= 16'h0000;
            14'h386c: oData <= 16'h0000;
            14'h386d: oData <= 16'h0000;
            14'h386e: oData <= 16'h0000;
            14'h386f: oData <= 16'h0000;
            14'h3870: oData <= 16'h0000;
            14'h3871: oData <= 16'h0000;
            14'h3872: oData <= 16'h0000;
            14'h3873: oData <= 16'h0000;
            14'h3874: oData <= 16'h0000;
            14'h3875: oData <= 16'h0000;
            14'h3876: oData <= 16'h0000;
            14'h3877: oData <= 16'h0000;
            14'h3878: oData <= 16'h0000;
            14'h3879: oData <= 16'h0000;
            14'h387a: oData <= 16'h0000;
            14'h387b: oData <= 16'h0000;
            14'h387c: oData <= 16'h0000;
            14'h387d: oData <= 16'h0000;
            14'h387e: oData <= 16'h0000;
            14'h387f: oData <= 16'h0000;
            14'h3880: oData <= 16'h0000;
            14'h3881: oData <= 16'h0000;
            14'h3882: oData <= 16'h0000;
            14'h3883: oData <= 16'h0000;
            14'h3884: oData <= 16'h0000;
            14'h3885: oData <= 16'h0000;
            14'h3886: oData <= 16'h0000;
            14'h3887: oData <= 16'h0000;
            14'h3888: oData <= 16'h0000;
            14'h3889: oData <= 16'h0000;
            14'h388a: oData <= 16'h0000;
            14'h388b: oData <= 16'h0000;
            14'h388c: oData <= 16'h0000;
            14'h388d: oData <= 16'h0000;
            14'h388e: oData <= 16'h0000;
            14'h388f: oData <= 16'h0000;
            14'h3890: oData <= 16'h0000;
            14'h3891: oData <= 16'h0000;
            14'h3892: oData <= 16'h0000;
            14'h3893: oData <= 16'h0000;
            14'h3894: oData <= 16'h0000;
            14'h3895: oData <= 16'h0000;
            14'h3896: oData <= 16'h0000;
            14'h3897: oData <= 16'h0000;
            14'h3898: oData <= 16'h0000;
            14'h3899: oData <= 16'h0000;
            14'h389a: oData <= 16'h0000;
            14'h389b: oData <= 16'h0000;
            14'h389c: oData <= 16'h0000;
            14'h389d: oData <= 16'h0000;
            14'h389e: oData <= 16'h0000;
            14'h389f: oData <= 16'h0000;
            14'h38a0: oData <= 16'h0000;
            14'h38a1: oData <= 16'h0000;
            14'h38a2: oData <= 16'h0000;
            14'h38a3: oData <= 16'h0000;
            14'h38a4: oData <= 16'h0000;
            14'h38a5: oData <= 16'h0000;
            14'h38a6: oData <= 16'h0000;
            14'h38a7: oData <= 16'h0000;
            14'h38a8: oData <= 16'h0000;
            14'h38a9: oData <= 16'h0000;
            14'h38aa: oData <= 16'h0000;
            14'h38ab: oData <= 16'h0000;
            14'h38ac: oData <= 16'h0000;
            14'h38ad: oData <= 16'h0000;
            14'h38ae: oData <= 16'h0000;
            14'h38af: oData <= 16'h0000;
            14'h38b0: oData <= 16'h0000;
            14'h38b1: oData <= 16'h0000;
            14'h38b2: oData <= 16'h0000;
            14'h38b3: oData <= 16'h0000;
            14'h38b4: oData <= 16'h0000;
            14'h38b5: oData <= 16'h0000;
            14'h38b6: oData <= 16'h0000;
            14'h38b7: oData <= 16'h0000;
            14'h38b8: oData <= 16'h0000;
            14'h38b9: oData <= 16'h0000;
            14'h38ba: oData <= 16'h0000;
            14'h38bb: oData <= 16'h0000;
            14'h38bc: oData <= 16'h0000;
            14'h38bd: oData <= 16'h0000;
            14'h38be: oData <= 16'h0000;
            14'h38bf: oData <= 16'h0000;
            14'h38c0: oData <= 16'h0000;
            14'h38c1: oData <= 16'h0000;
            14'h38c2: oData <= 16'h0000;
            14'h38c3: oData <= 16'h0000;
            14'h38c4: oData <= 16'h0000;
            14'h38c5: oData <= 16'h0000;
            14'h38c6: oData <= 16'h0000;
            14'h38c7: oData <= 16'h0000;
            14'h38c8: oData <= 16'h0000;
            14'h38c9: oData <= 16'h0000;
            14'h38ca: oData <= 16'h0000;
            14'h38cb: oData <= 16'h0000;
            14'h38cc: oData <= 16'h0000;
            14'h38cd: oData <= 16'h0000;
            14'h38ce: oData <= 16'h0000;
            14'h38cf: oData <= 16'h0000;
            14'h38d0: oData <= 16'h0000;
            14'h38d1: oData <= 16'h0000;
            14'h38d2: oData <= 16'h0000;
            14'h38d3: oData <= 16'h0000;
            14'h38d4: oData <= 16'h0000;
            14'h38d5: oData <= 16'h0000;
            14'h38d6: oData <= 16'h0000;
            14'h38d7: oData <= 16'h0000;
            14'h38d8: oData <= 16'h0000;
            14'h38d9: oData <= 16'h0000;
            14'h38da: oData <= 16'h0000;
            14'h38db: oData <= 16'h0000;
            14'h38dc: oData <= 16'h0000;
            14'h38dd: oData <= 16'h0000;
            14'h38de: oData <= 16'h0000;
            14'h38df: oData <= 16'h0000;
            14'h38e0: oData <= 16'h0000;
            14'h38e1: oData <= 16'h0000;
            14'h38e2: oData <= 16'h0000;
            14'h38e3: oData <= 16'h0000;
            14'h38e4: oData <= 16'h0000;
            14'h38e5: oData <= 16'h0000;
            14'h38e6: oData <= 16'h0000;
            14'h38e7: oData <= 16'h0000;
            14'h38e8: oData <= 16'h0000;
            14'h38e9: oData <= 16'h0000;
            14'h38ea: oData <= 16'h0000;
            14'h38eb: oData <= 16'h0000;
            14'h38ec: oData <= 16'h0000;
            14'h38ed: oData <= 16'h0000;
            14'h38ee: oData <= 16'h0000;
            14'h38ef: oData <= 16'h0000;
            14'h38f0: oData <= 16'h0000;
            14'h38f1: oData <= 16'h0000;
            14'h38f2: oData <= 16'h0000;
            14'h38f3: oData <= 16'h0000;
            14'h38f4: oData <= 16'h0000;
            14'h38f5: oData <= 16'h0000;
            14'h38f6: oData <= 16'h0000;
            14'h38f7: oData <= 16'h0000;
            14'h38f8: oData <= 16'h0000;
            14'h38f9: oData <= 16'h0000;
            14'h38fa: oData <= 16'h0000;
            14'h38fb: oData <= 16'h0000;
            14'h38fc: oData <= 16'h0000;
            14'h38fd: oData <= 16'h0000;
            14'h38fe: oData <= 16'h0000;
            14'h38ff: oData <= 16'h0000;
            14'h3900: oData <= 16'h0000;
            14'h3901: oData <= 16'h0000;
            14'h3902: oData <= 16'h0000;
            14'h3903: oData <= 16'h0000;
            14'h3904: oData <= 16'h0000;
            14'h3905: oData <= 16'h0000;
            14'h3906: oData <= 16'h0000;
            14'h3907: oData <= 16'h0000;
            14'h3908: oData <= 16'h0000;
            14'h3909: oData <= 16'h0000;
            14'h390a: oData <= 16'h0000;
            14'h390b: oData <= 16'h0000;
            14'h390c: oData <= 16'h0000;
            14'h390d: oData <= 16'h0000;
            14'h390e: oData <= 16'h0000;
            14'h390f: oData <= 16'h0000;
            14'h3910: oData <= 16'h0000;
            14'h3911: oData <= 16'h0000;
            14'h3912: oData <= 16'h0000;
            14'h3913: oData <= 16'h0000;
            14'h3914: oData <= 16'h0000;
            14'h3915: oData <= 16'h0000;
            14'h3916: oData <= 16'h0000;
            14'h3917: oData <= 16'h0000;
            14'h3918: oData <= 16'h0000;
            14'h3919: oData <= 16'h0000;
            14'h391a: oData <= 16'h0000;
            14'h391b: oData <= 16'h0000;
            14'h391c: oData <= 16'h0000;
            14'h391d: oData <= 16'h0000;
            14'h391e: oData <= 16'h0000;
            14'h391f: oData <= 16'h0000;
            14'h3920: oData <= 16'h0000;
            14'h3921: oData <= 16'h0000;
            14'h3922: oData <= 16'h0000;
            14'h3923: oData <= 16'h0000;
            14'h3924: oData <= 16'h0000;
            14'h3925: oData <= 16'h0000;
            14'h3926: oData <= 16'h0000;
            14'h3927: oData <= 16'h0000;
            14'h3928: oData <= 16'h0000;
            14'h3929: oData <= 16'h0000;
            14'h392a: oData <= 16'h0000;
            14'h392b: oData <= 16'h0000;
            14'h392c: oData <= 16'h0000;
            14'h392d: oData <= 16'h0000;
            14'h392e: oData <= 16'h0000;
            14'h392f: oData <= 16'h0000;
            14'h3930: oData <= 16'h0000;
            14'h3931: oData <= 16'h0000;
            14'h3932: oData <= 16'h0000;
            14'h3933: oData <= 16'h0000;
            14'h3934: oData <= 16'h0000;
            14'h3935: oData <= 16'h0000;
            14'h3936: oData <= 16'h0000;
            14'h3937: oData <= 16'h0000;
            14'h3938: oData <= 16'h0000;
            14'h3939: oData <= 16'h0000;
            14'h393a: oData <= 16'h0000;
            14'h393b: oData <= 16'h0000;
            14'h393c: oData <= 16'h0000;
            14'h393d: oData <= 16'h0000;
            14'h393e: oData <= 16'h0000;
            14'h393f: oData <= 16'h0000;
            14'h3940: oData <= 16'h0000;
            14'h3941: oData <= 16'h0000;
            14'h3942: oData <= 16'h0000;
            14'h3943: oData <= 16'h0000;
            14'h3944: oData <= 16'h0000;
            14'h3945: oData <= 16'h0000;
            14'h3946: oData <= 16'h0000;
            14'h3947: oData <= 16'h0000;
            14'h3948: oData <= 16'h0000;
            14'h3949: oData <= 16'h0000;
            14'h394a: oData <= 16'h0000;
            14'h394b: oData <= 16'h0000;
            14'h394c: oData <= 16'h0000;
            14'h394d: oData <= 16'h0000;
            14'h394e: oData <= 16'h0000;
            14'h394f: oData <= 16'h0000;
            14'h3950: oData <= 16'h0000;
            14'h3951: oData <= 16'h0000;
            14'h3952: oData <= 16'h0000;
            14'h3953: oData <= 16'h0000;
            14'h3954: oData <= 16'h0000;
            14'h3955: oData <= 16'h0000;
            14'h3956: oData <= 16'h0000;
            14'h3957: oData <= 16'h0000;
            14'h3958: oData <= 16'h0000;
            14'h3959: oData <= 16'h0000;
            14'h395a: oData <= 16'h0000;
            14'h395b: oData <= 16'h0000;
            14'h395c: oData <= 16'h0000;
            14'h395d: oData <= 16'h0000;
            14'h395e: oData <= 16'h0000;
            14'h395f: oData <= 16'h0000;
            14'h3960: oData <= 16'h0000;
            14'h3961: oData <= 16'h0000;
            14'h3962: oData <= 16'h0000;
            14'h3963: oData <= 16'h0000;
            14'h3964: oData <= 16'h0000;
            14'h3965: oData <= 16'h0000;
            14'h3966: oData <= 16'h0000;
            14'h3967: oData <= 16'h0000;
            14'h3968: oData <= 16'h0000;
            14'h3969: oData <= 16'h0000;
            14'h396a: oData <= 16'h0000;
            14'h396b: oData <= 16'h0000;
            14'h396c: oData <= 16'h0000;
            14'h396d: oData <= 16'h0000;
            14'h396e: oData <= 16'h0000;
            14'h396f: oData <= 16'h0000;
            14'h3970: oData <= 16'h0000;
            14'h3971: oData <= 16'h0000;
            14'h3972: oData <= 16'h0000;
            14'h3973: oData <= 16'h0000;
            14'h3974: oData <= 16'h0000;
            14'h3975: oData <= 16'h0000;
            14'h3976: oData <= 16'h0000;
            14'h3977: oData <= 16'h0000;
            14'h3978: oData <= 16'h0000;
            14'h3979: oData <= 16'h0000;
            14'h397a: oData <= 16'h0000;
            14'h397b: oData <= 16'h0000;
            14'h397c: oData <= 16'h0000;
            14'h397d: oData <= 16'h0000;
            14'h397e: oData <= 16'h0000;
            14'h397f: oData <= 16'h0000;
            14'h3980: oData <= 16'h0000;
            14'h3981: oData <= 16'h0000;
            14'h3982: oData <= 16'h0000;
            14'h3983: oData <= 16'h0000;
            14'h3984: oData <= 16'h0000;
            14'h3985: oData <= 16'h0000;
            14'h3986: oData <= 16'h0000;
            14'h3987: oData <= 16'h0000;
            14'h3988: oData <= 16'h0000;
            14'h3989: oData <= 16'h0000;
            14'h398a: oData <= 16'h0000;
            14'h398b: oData <= 16'h0000;
            14'h398c: oData <= 16'h0000;
            14'h398d: oData <= 16'h0000;
            14'h398e: oData <= 16'h0000;
            14'h398f: oData <= 16'h0000;
            14'h3990: oData <= 16'h0000;
            14'h3991: oData <= 16'h0000;
            14'h3992: oData <= 16'h0000;
            14'h3993: oData <= 16'h0000;
            14'h3994: oData <= 16'h0000;
            14'h3995: oData <= 16'h0000;
            14'h3996: oData <= 16'h0000;
            14'h3997: oData <= 16'h0000;
            14'h3998: oData <= 16'h0000;
            14'h3999: oData <= 16'h0000;
            14'h399a: oData <= 16'h0000;
            14'h399b: oData <= 16'h0000;
            14'h399c: oData <= 16'h0000;
            14'h399d: oData <= 16'h0000;
            14'h399e: oData <= 16'h0000;
            14'h399f: oData <= 16'h0000;
            14'h39a0: oData <= 16'h0000;
            14'h39a1: oData <= 16'h0000;
            14'h39a2: oData <= 16'h0000;
            14'h39a3: oData <= 16'h0000;
            14'h39a4: oData <= 16'h0000;
            14'h39a5: oData <= 16'h0000;
            14'h39a6: oData <= 16'h0000;
            14'h39a7: oData <= 16'h0000;
            14'h39a8: oData <= 16'h0000;
            14'h39a9: oData <= 16'h0000;
            14'h39aa: oData <= 16'h0000;
            14'h39ab: oData <= 16'h0000;
            14'h39ac: oData <= 16'h0000;
            14'h39ad: oData <= 16'h0000;
            14'h39ae: oData <= 16'h0000;
            14'h39af: oData <= 16'h0000;
            14'h39b0: oData <= 16'h0000;
            14'h39b1: oData <= 16'h0000;
            14'h39b2: oData <= 16'h0000;
            14'h39b3: oData <= 16'h0000;
            14'h39b4: oData <= 16'h0000;
            14'h39b5: oData <= 16'h0000;
            14'h39b6: oData <= 16'h0000;
            14'h39b7: oData <= 16'h0000;
            14'h39b8: oData <= 16'h0000;
            14'h39b9: oData <= 16'h0000;
            14'h39ba: oData <= 16'h0000;
            14'h39bb: oData <= 16'h0000;
            14'h39bc: oData <= 16'h0000;
            14'h39bd: oData <= 16'h0000;
            14'h39be: oData <= 16'h0000;
            14'h39bf: oData <= 16'h0000;
            14'h39c0: oData <= 16'h0000;
            14'h39c1: oData <= 16'h0000;
            14'h39c2: oData <= 16'h0000;
            14'h39c3: oData <= 16'h0000;
            14'h39c4: oData <= 16'h0000;
            14'h39c5: oData <= 16'h0000;
            14'h39c6: oData <= 16'h0000;
            14'h39c7: oData <= 16'h0000;
            14'h39c8: oData <= 16'h0000;
            14'h39c9: oData <= 16'h0000;
            14'h39ca: oData <= 16'h0000;
            14'h39cb: oData <= 16'h0000;
            14'h39cc: oData <= 16'h0000;
            14'h39cd: oData <= 16'h0000;
            14'h39ce: oData <= 16'h0000;
            14'h39cf: oData <= 16'h0000;
            14'h39d0: oData <= 16'h0000;
            14'h39d1: oData <= 16'h0000;
            14'h39d2: oData <= 16'h0000;
            14'h39d3: oData <= 16'h0000;
            14'h39d4: oData <= 16'h0000;
            14'h39d5: oData <= 16'h0000;
            14'h39d6: oData <= 16'h0000;
            14'h39d7: oData <= 16'h0000;
            14'h39d8: oData <= 16'h0000;
            14'h39d9: oData <= 16'h0000;
            14'h39da: oData <= 16'h0000;
            14'h39db: oData <= 16'h0000;
            14'h39dc: oData <= 16'h0000;
            14'h39dd: oData <= 16'h0000;
            14'h39de: oData <= 16'h0000;
            14'h39df: oData <= 16'h0000;
            14'h39e0: oData <= 16'h0000;
            14'h39e1: oData <= 16'h0000;
            14'h39e2: oData <= 16'h0000;
            14'h39e3: oData <= 16'h0000;
            14'h39e4: oData <= 16'h0000;
            14'h39e5: oData <= 16'h0000;
            14'h39e6: oData <= 16'h0000;
            14'h39e7: oData <= 16'h0000;
            14'h39e8: oData <= 16'h0000;
            14'h39e9: oData <= 16'h0000;
            14'h39ea: oData <= 16'h0000;
            14'h39eb: oData <= 16'h0000;
            14'h39ec: oData <= 16'h0000;
            14'h39ed: oData <= 16'h0000;
            14'h39ee: oData <= 16'h0000;
            14'h39ef: oData <= 16'h0000;
            14'h39f0: oData <= 16'h0000;
            14'h39f1: oData <= 16'h0000;
            14'h39f2: oData <= 16'h0000;
            14'h39f3: oData <= 16'h0000;
            14'h39f4: oData <= 16'h0000;
            14'h39f5: oData <= 16'h0000;
            14'h39f6: oData <= 16'h0000;
            14'h39f7: oData <= 16'h0000;
            14'h39f8: oData <= 16'h0000;
            14'h39f9: oData <= 16'h0000;
            14'h39fa: oData <= 16'h0000;
            14'h39fb: oData <= 16'h0000;
            14'h39fc: oData <= 16'h0000;
            14'h39fd: oData <= 16'h0000;
            14'h39fe: oData <= 16'h0000;
            14'h39ff: oData <= 16'h0000;
            14'h3a00: oData <= 16'h0000;
            14'h3a01: oData <= 16'h0000;
            14'h3a02: oData <= 16'h0000;
            14'h3a03: oData <= 16'h0000;
            14'h3a04: oData <= 16'h0000;
            14'h3a05: oData <= 16'h0000;
            14'h3a06: oData <= 16'h0000;
            14'h3a07: oData <= 16'h0000;
            14'h3a08: oData <= 16'h0000;
            14'h3a09: oData <= 16'h0000;
            14'h3a0a: oData <= 16'h0000;
            14'h3a0b: oData <= 16'h0000;
            14'h3a0c: oData <= 16'h0000;
            14'h3a0d: oData <= 16'h0000;
            14'h3a0e: oData <= 16'h0000;
            14'h3a0f: oData <= 16'h0000;
            14'h3a10: oData <= 16'h0000;
            14'h3a11: oData <= 16'h0000;
            14'h3a12: oData <= 16'h0000;
            14'h3a13: oData <= 16'h0000;
            14'h3a14: oData <= 16'h0000;
            14'h3a15: oData <= 16'h0000;
            14'h3a16: oData <= 16'h0000;
            14'h3a17: oData <= 16'h0000;
            14'h3a18: oData <= 16'h0000;
            14'h3a19: oData <= 16'h0000;
            14'h3a1a: oData <= 16'h0000;
            14'h3a1b: oData <= 16'h0000;
            14'h3a1c: oData <= 16'h0000;
            14'h3a1d: oData <= 16'h0000;
            14'h3a1e: oData <= 16'h0000;
            14'h3a1f: oData <= 16'h0000;
            14'h3a20: oData <= 16'h0000;
            14'h3a21: oData <= 16'h0000;
            14'h3a22: oData <= 16'h0000;
            14'h3a23: oData <= 16'h0000;
            14'h3a24: oData <= 16'h0000;
            14'h3a25: oData <= 16'h0000;
            14'h3a26: oData <= 16'h0000;
            14'h3a27: oData <= 16'h0000;
            14'h3a28: oData <= 16'h0000;
            14'h3a29: oData <= 16'h0000;
            14'h3a2a: oData <= 16'h0000;
            14'h3a2b: oData <= 16'h0000;
            14'h3a2c: oData <= 16'h0000;
            14'h3a2d: oData <= 16'h0000;
            14'h3a2e: oData <= 16'h0000;
            14'h3a2f: oData <= 16'h0000;
            14'h3a30: oData <= 16'h0000;
            14'h3a31: oData <= 16'h0000;
            14'h3a32: oData <= 16'h0000;
            14'h3a33: oData <= 16'h0000;
            14'h3a34: oData <= 16'h0000;
            14'h3a35: oData <= 16'h0000;
            14'h3a36: oData <= 16'h0000;
            14'h3a37: oData <= 16'h0000;
            14'h3a38: oData <= 16'h0000;
            14'h3a39: oData <= 16'h0000;
            14'h3a3a: oData <= 16'h0000;
            14'h3a3b: oData <= 16'h0000;
            14'h3a3c: oData <= 16'h0000;
            14'h3a3d: oData <= 16'h0000;
            14'h3a3e: oData <= 16'h0000;
            14'h3a3f: oData <= 16'h0000;
            14'h3a40: oData <= 16'h0000;
            14'h3a41: oData <= 16'h0000;
            14'h3a42: oData <= 16'h0000;
            14'h3a43: oData <= 16'h0000;
            14'h3a44: oData <= 16'h0000;
            14'h3a45: oData <= 16'h0000;
            14'h3a46: oData <= 16'h0000;
            14'h3a47: oData <= 16'h0000;
            14'h3a48: oData <= 16'h0000;
            14'h3a49: oData <= 16'h0000;
            14'h3a4a: oData <= 16'h0000;
            14'h3a4b: oData <= 16'h0000;
            14'h3a4c: oData <= 16'h0000;
            14'h3a4d: oData <= 16'h0000;
            14'h3a4e: oData <= 16'h0000;
            14'h3a4f: oData <= 16'h0000;
            14'h3a50: oData <= 16'h0000;
            14'h3a51: oData <= 16'h0000;
            14'h3a52: oData <= 16'h0000;
            14'h3a53: oData <= 16'h0000;
            14'h3a54: oData <= 16'h0000;
            14'h3a55: oData <= 16'h0000;
            14'h3a56: oData <= 16'h0000;
            14'h3a57: oData <= 16'h0000;
            14'h3a58: oData <= 16'h0000;
            14'h3a59: oData <= 16'h0000;
            14'h3a5a: oData <= 16'h0000;
            14'h3a5b: oData <= 16'h0000;
            14'h3a5c: oData <= 16'h0000;
            14'h3a5d: oData <= 16'h0000;
            14'h3a5e: oData <= 16'h0000;
            14'h3a5f: oData <= 16'h0000;
            14'h3a60: oData <= 16'h0000;
            14'h3a61: oData <= 16'h0000;
            14'h3a62: oData <= 16'h0000;
            14'h3a63: oData <= 16'h0000;
            14'h3a64: oData <= 16'h0000;
            14'h3a65: oData <= 16'h0000;
            14'h3a66: oData <= 16'h0000;
            14'h3a67: oData <= 16'h0000;
            14'h3a68: oData <= 16'h0000;
            14'h3a69: oData <= 16'h0000;
            14'h3a6a: oData <= 16'h0000;
            14'h3a6b: oData <= 16'h0000;
            14'h3a6c: oData <= 16'h0000;
            14'h3a6d: oData <= 16'h0000;
            14'h3a6e: oData <= 16'h0000;
            14'h3a6f: oData <= 16'h0000;
            14'h3a70: oData <= 16'h0000;
            14'h3a71: oData <= 16'h0000;
            14'h3a72: oData <= 16'h0000;
            14'h3a73: oData <= 16'h0000;
            14'h3a74: oData <= 16'h0000;
            14'h3a75: oData <= 16'h0000;
            14'h3a76: oData <= 16'h0000;
            14'h3a77: oData <= 16'h0000;
            14'h3a78: oData <= 16'h0000;
            14'h3a79: oData <= 16'h0000;
            14'h3a7a: oData <= 16'h0000;
            14'h3a7b: oData <= 16'h0000;
            14'h3a7c: oData <= 16'h0000;
            14'h3a7d: oData <= 16'h0000;
            14'h3a7e: oData <= 16'h0000;
            14'h3a7f: oData <= 16'h0000;
            14'h3a80: oData <= 16'h0000;
            14'h3a81: oData <= 16'h0000;
            14'h3a82: oData <= 16'h0000;
            14'h3a83: oData <= 16'h0000;
            14'h3a84: oData <= 16'h0000;
            14'h3a85: oData <= 16'h0000;
            14'h3a86: oData <= 16'h0000;
            14'h3a87: oData <= 16'h0000;
            14'h3a88: oData <= 16'h0000;
            14'h3a89: oData <= 16'h0000;
            14'h3a8a: oData <= 16'h0000;
            14'h3a8b: oData <= 16'h0000;
            14'h3a8c: oData <= 16'h0000;
            14'h3a8d: oData <= 16'h0000;
            14'h3a8e: oData <= 16'h0000;
            14'h3a8f: oData <= 16'h0000;
            14'h3a90: oData <= 16'h0000;
            14'h3a91: oData <= 16'h0000;
            14'h3a92: oData <= 16'h0000;
            14'h3a93: oData <= 16'h0000;
            14'h3a94: oData <= 16'h0000;
            14'h3a95: oData <= 16'h0000;
            14'h3a96: oData <= 16'h0000;
            14'h3a97: oData <= 16'h0000;
            14'h3a98: oData <= 16'h0000;
            14'h3a99: oData <= 16'h0000;
            14'h3a9a: oData <= 16'h0000;
            14'h3a9b: oData <= 16'h0000;
            14'h3a9c: oData <= 16'h0000;
            14'h3a9d: oData <= 16'h0000;
            14'h3a9e: oData <= 16'h0000;
            14'h3a9f: oData <= 16'h0000;
            14'h3aa0: oData <= 16'h0000;
            14'h3aa1: oData <= 16'h0000;
            14'h3aa2: oData <= 16'h0000;
            14'h3aa3: oData <= 16'h0000;
            14'h3aa4: oData <= 16'h0000;
            14'h3aa5: oData <= 16'h0000;
            14'h3aa6: oData <= 16'h0000;
            14'h3aa7: oData <= 16'h0000;
            14'h3aa8: oData <= 16'h0000;
            14'h3aa9: oData <= 16'h0000;
            14'h3aaa: oData <= 16'h0000;
            14'h3aab: oData <= 16'h0000;
            14'h3aac: oData <= 16'h0000;
            14'h3aad: oData <= 16'h0000;
            14'h3aae: oData <= 16'h0000;
            14'h3aaf: oData <= 16'h0000;
            14'h3ab0: oData <= 16'h0000;
            14'h3ab1: oData <= 16'h0000;
            14'h3ab2: oData <= 16'h0000;
            14'h3ab3: oData <= 16'h0000;
            14'h3ab4: oData <= 16'h0000;
            14'h3ab5: oData <= 16'h0000;
            14'h3ab6: oData <= 16'h0000;
            14'h3ab7: oData <= 16'h0000;
            14'h3ab8: oData <= 16'h0000;
            14'h3ab9: oData <= 16'h0000;
            14'h3aba: oData <= 16'h0000;
            14'h3abb: oData <= 16'h0000;
            14'h3abc: oData <= 16'h0000;
            14'h3abd: oData <= 16'h0000;
            14'h3abe: oData <= 16'h0000;
            14'h3abf: oData <= 16'h0000;
            14'h3ac0: oData <= 16'h0000;
            14'h3ac1: oData <= 16'h0000;
            14'h3ac2: oData <= 16'h0000;
            14'h3ac3: oData <= 16'h0000;
            14'h3ac4: oData <= 16'h0000;
            14'h3ac5: oData <= 16'h0000;
            14'h3ac6: oData <= 16'h0000;
            14'h3ac7: oData <= 16'h0000;
            14'h3ac8: oData <= 16'h0000;
            14'h3ac9: oData <= 16'h0000;
            14'h3aca: oData <= 16'h0000;
            14'h3acb: oData <= 16'h0000;
            14'h3acc: oData <= 16'h0000;
            14'h3acd: oData <= 16'h0000;
            14'h3ace: oData <= 16'h0000;
            14'h3acf: oData <= 16'h0000;
            14'h3ad0: oData <= 16'h0000;
            14'h3ad1: oData <= 16'h0000;
            14'h3ad2: oData <= 16'h0000;
            14'h3ad3: oData <= 16'h0000;
            14'h3ad4: oData <= 16'h0000;
            14'h3ad5: oData <= 16'h0000;
            14'h3ad6: oData <= 16'h0000;
            14'h3ad7: oData <= 16'h0000;
            14'h3ad8: oData <= 16'h0000;
            14'h3ad9: oData <= 16'h0000;
            14'h3ada: oData <= 16'h0000;
            14'h3adb: oData <= 16'h0000;
            14'h3adc: oData <= 16'h0000;
            14'h3add: oData <= 16'h0000;
            14'h3ade: oData <= 16'h0000;
            14'h3adf: oData <= 16'h0000;
            14'h3ae0: oData <= 16'h0000;
            14'h3ae1: oData <= 16'h0000;
            14'h3ae2: oData <= 16'h0000;
            14'h3ae3: oData <= 16'h0000;
            14'h3ae4: oData <= 16'h0000;
            14'h3ae5: oData <= 16'h0000;
            14'h3ae6: oData <= 16'h0000;
            14'h3ae7: oData <= 16'h0000;
            14'h3ae8: oData <= 16'h0000;
            14'h3ae9: oData <= 16'h0000;
            14'h3aea: oData <= 16'h0000;
            14'h3aeb: oData <= 16'h0000;
            14'h3aec: oData <= 16'h0000;
            14'h3aed: oData <= 16'h0000;
            14'h3aee: oData <= 16'h0000;
            14'h3aef: oData <= 16'h0000;
            14'h3af0: oData <= 16'h0000;
            14'h3af1: oData <= 16'h0000;
            14'h3af2: oData <= 16'h0000;
            14'h3af3: oData <= 16'h0000;
            14'h3af4: oData <= 16'h0000;
            14'h3af5: oData <= 16'h0000;
            14'h3af6: oData <= 16'h0000;
            14'h3af7: oData <= 16'h0000;
            14'h3af8: oData <= 16'h0000;
            14'h3af9: oData <= 16'h0000;
            14'h3afa: oData <= 16'h0000;
            14'h3afb: oData <= 16'h0000;
            14'h3afc: oData <= 16'h0000;
            14'h3afd: oData <= 16'h0000;
            14'h3afe: oData <= 16'h0000;
            14'h3aff: oData <= 16'h0000;
            14'h3b00: oData <= 16'h0000;
            14'h3b01: oData <= 16'h0000;
            14'h3b02: oData <= 16'h0000;
            14'h3b03: oData <= 16'h0000;
            14'h3b04: oData <= 16'h0000;
            14'h3b05: oData <= 16'h0000;
            14'h3b06: oData <= 16'h0000;
            14'h3b07: oData <= 16'h0000;
            14'h3b08: oData <= 16'h0000;
            14'h3b09: oData <= 16'h0000;
            14'h3b0a: oData <= 16'h0000;
            14'h3b0b: oData <= 16'h0000;
            14'h3b0c: oData <= 16'h0000;
            14'h3b0d: oData <= 16'h0000;
            14'h3b0e: oData <= 16'h0000;
            14'h3b0f: oData <= 16'h0000;
            14'h3b10: oData <= 16'h0000;
            14'h3b11: oData <= 16'h0000;
            14'h3b12: oData <= 16'h0000;
            14'h3b13: oData <= 16'h0000;
            14'h3b14: oData <= 16'h0000;
            14'h3b15: oData <= 16'h0000;
            14'h3b16: oData <= 16'h0000;
            14'h3b17: oData <= 16'h0000;
            14'h3b18: oData <= 16'h0000;
            14'h3b19: oData <= 16'h0000;
            14'h3b1a: oData <= 16'h0000;
            14'h3b1b: oData <= 16'h0000;
            14'h3b1c: oData <= 16'h0000;
            14'h3b1d: oData <= 16'h0000;
            14'h3b1e: oData <= 16'h0000;
            14'h3b1f: oData <= 16'h0000;
            14'h3b20: oData <= 16'h0000;
            14'h3b21: oData <= 16'h0000;
            14'h3b22: oData <= 16'h0000;
            14'h3b23: oData <= 16'h0000;
            14'h3b24: oData <= 16'h0000;
            14'h3b25: oData <= 16'h0000;
            14'h3b26: oData <= 16'h0000;
            14'h3b27: oData <= 16'h0000;
            14'h3b28: oData <= 16'h0000;
            14'h3b29: oData <= 16'h0000;
            14'h3b2a: oData <= 16'h0000;
            14'h3b2b: oData <= 16'h0000;
            14'h3b2c: oData <= 16'h0000;
            14'h3b2d: oData <= 16'h0000;
            14'h3b2e: oData <= 16'h0000;
            14'h3b2f: oData <= 16'h0000;
            14'h3b30: oData <= 16'h0000;
            14'h3b31: oData <= 16'h0000;
            14'h3b32: oData <= 16'h0000;
            14'h3b33: oData <= 16'h0000;
            14'h3b34: oData <= 16'h0000;
            14'h3b35: oData <= 16'h0000;
            14'h3b36: oData <= 16'h0000;
            14'h3b37: oData <= 16'h0000;
            14'h3b38: oData <= 16'h0000;
            14'h3b39: oData <= 16'h0000;
            14'h3b3a: oData <= 16'h0000;
            14'h3b3b: oData <= 16'h0000;
            14'h3b3c: oData <= 16'h0000;
            14'h3b3d: oData <= 16'h0000;
            14'h3b3e: oData <= 16'h0000;
            14'h3b3f: oData <= 16'h0000;
            14'h3b40: oData <= 16'h0000;
            14'h3b41: oData <= 16'h0000;
            14'h3b42: oData <= 16'h0000;
            14'h3b43: oData <= 16'h0000;
            14'h3b44: oData <= 16'h0000;
            14'h3b45: oData <= 16'h0000;
            14'h3b46: oData <= 16'h0000;
            14'h3b47: oData <= 16'h0000;
            14'h3b48: oData <= 16'h0000;
            14'h3b49: oData <= 16'h0000;
            14'h3b4a: oData <= 16'h0000;
            14'h3b4b: oData <= 16'h0000;
            14'h3b4c: oData <= 16'h0000;
            14'h3b4d: oData <= 16'h0000;
            14'h3b4e: oData <= 16'h0000;
            14'h3b4f: oData <= 16'h0000;
            14'h3b50: oData <= 16'h0000;
            14'h3b51: oData <= 16'h0000;
            14'h3b52: oData <= 16'h0000;
            14'h3b53: oData <= 16'h0000;
            14'h3b54: oData <= 16'h0000;
            14'h3b55: oData <= 16'h0000;
            14'h3b56: oData <= 16'h0000;
            14'h3b57: oData <= 16'h0000;
            14'h3b58: oData <= 16'h0000;
            14'h3b59: oData <= 16'h0000;
            14'h3b5a: oData <= 16'h0000;
            14'h3b5b: oData <= 16'h0000;
            14'h3b5c: oData <= 16'h0000;
            14'h3b5d: oData <= 16'h0000;
            14'h3b5e: oData <= 16'h0000;
            14'h3b5f: oData <= 16'h0000;
            14'h3b60: oData <= 16'h0000;
            14'h3b61: oData <= 16'h0000;
            14'h3b62: oData <= 16'h0000;
            14'h3b63: oData <= 16'h0000;
            14'h3b64: oData <= 16'h0000;
            14'h3b65: oData <= 16'h0000;
            14'h3b66: oData <= 16'h0000;
            14'h3b67: oData <= 16'h0000;
            14'h3b68: oData <= 16'h0000;
            14'h3b69: oData <= 16'h0000;
            14'h3b6a: oData <= 16'h0000;
            14'h3b6b: oData <= 16'h0000;
            14'h3b6c: oData <= 16'h0000;
            14'h3b6d: oData <= 16'h0000;
            14'h3b6e: oData <= 16'h0000;
            14'h3b6f: oData <= 16'h0000;
            14'h3b70: oData <= 16'h0000;
            14'h3b71: oData <= 16'h0000;
            14'h3b72: oData <= 16'h0000;
            14'h3b73: oData <= 16'h0000;
            14'h3b74: oData <= 16'h0000;
            14'h3b75: oData <= 16'h0000;
            14'h3b76: oData <= 16'h0000;
            14'h3b77: oData <= 16'h0000;
            14'h3b78: oData <= 16'h0000;
            14'h3b79: oData <= 16'h0000;
            14'h3b7a: oData <= 16'h0000;
            14'h3b7b: oData <= 16'h0000;
            14'h3b7c: oData <= 16'h0000;
            14'h3b7d: oData <= 16'h0000;
            14'h3b7e: oData <= 16'h0000;
            14'h3b7f: oData <= 16'h0000;
            14'h3b80: oData <= 16'h0000;
            14'h3b81: oData <= 16'h0000;
            14'h3b82: oData <= 16'h0000;
            14'h3b83: oData <= 16'h0000;
            14'h3b84: oData <= 16'h0000;
            14'h3b85: oData <= 16'h0000;
            14'h3b86: oData <= 16'h0000;
            14'h3b87: oData <= 16'h0000;
            14'h3b88: oData <= 16'h0000;
            14'h3b89: oData <= 16'h0000;
            14'h3b8a: oData <= 16'h0000;
            14'h3b8b: oData <= 16'h0000;
            14'h3b8c: oData <= 16'h0000;
            14'h3b8d: oData <= 16'h0000;
            14'h3b8e: oData <= 16'h0000;
            14'h3b8f: oData <= 16'h0000;
            14'h3b90: oData <= 16'h0000;
            14'h3b91: oData <= 16'h0000;
            14'h3b92: oData <= 16'h0000;
            14'h3b93: oData <= 16'h0000;
            14'h3b94: oData <= 16'h0000;
            14'h3b95: oData <= 16'h0000;
            14'h3b96: oData <= 16'h0000;
            14'h3b97: oData <= 16'h0000;
            14'h3b98: oData <= 16'h0000;
            14'h3b99: oData <= 16'h0000;
            14'h3b9a: oData <= 16'h0000;
            14'h3b9b: oData <= 16'h0000;
            14'h3b9c: oData <= 16'h0000;
            14'h3b9d: oData <= 16'h0000;
            14'h3b9e: oData <= 16'h0000;
            14'h3b9f: oData <= 16'h0000;
            14'h3ba0: oData <= 16'h0000;
            14'h3ba1: oData <= 16'h0000;
            14'h3ba2: oData <= 16'h0000;
            14'h3ba3: oData <= 16'h0000;
            14'h3ba4: oData <= 16'h0000;
            14'h3ba5: oData <= 16'h0000;
            14'h3ba6: oData <= 16'h0000;
            14'h3ba7: oData <= 16'h0000;
            14'h3ba8: oData <= 16'h0000;
            14'h3ba9: oData <= 16'h0000;
            14'h3baa: oData <= 16'h0000;
            14'h3bab: oData <= 16'h0000;
            14'h3bac: oData <= 16'h0000;
            14'h3bad: oData <= 16'h0000;
            14'h3bae: oData <= 16'h0000;
            14'h3baf: oData <= 16'h0000;
            14'h3bb0: oData <= 16'h0000;
            14'h3bb1: oData <= 16'h0000;
            14'h3bb2: oData <= 16'h0000;
            14'h3bb3: oData <= 16'h0000;
            14'h3bb4: oData <= 16'h0000;
            14'h3bb5: oData <= 16'h0000;
            14'h3bb6: oData <= 16'h0000;
            14'h3bb7: oData <= 16'h0000;
            14'h3bb8: oData <= 16'h0000;
            14'h3bb9: oData <= 16'h0000;
            14'h3bba: oData <= 16'h0000;
            14'h3bbb: oData <= 16'h0000;
            14'h3bbc: oData <= 16'h0000;
            14'h3bbd: oData <= 16'h0000;
            14'h3bbe: oData <= 16'h0000;
            14'h3bbf: oData <= 16'h0000;
            14'h3bc0: oData <= 16'h0000;
            14'h3bc1: oData <= 16'h0000;
            14'h3bc2: oData <= 16'h0000;
            14'h3bc3: oData <= 16'h0000;
            14'h3bc4: oData <= 16'h0000;
            14'h3bc5: oData <= 16'h0000;
            14'h3bc6: oData <= 16'h0000;
            14'h3bc7: oData <= 16'h0000;
            14'h3bc8: oData <= 16'h0000;
            14'h3bc9: oData <= 16'h0000;
            14'h3bca: oData <= 16'h0000;
            14'h3bcb: oData <= 16'h0000;
            14'h3bcc: oData <= 16'h0000;
            14'h3bcd: oData <= 16'h0000;
            14'h3bce: oData <= 16'h0000;
            14'h3bcf: oData <= 16'h0000;
            14'h3bd0: oData <= 16'h0000;
            14'h3bd1: oData <= 16'h0000;
            14'h3bd2: oData <= 16'h0000;
            14'h3bd3: oData <= 16'h0000;
            14'h3bd4: oData <= 16'h0000;
            14'h3bd5: oData <= 16'h0000;
            14'h3bd6: oData <= 16'h0000;
            14'h3bd7: oData <= 16'h0000;
            14'h3bd8: oData <= 16'h0000;
            14'h3bd9: oData <= 16'h0000;
            14'h3bda: oData <= 16'h0000;
            14'h3bdb: oData <= 16'h0000;
            14'h3bdc: oData <= 16'h0000;
            14'h3bdd: oData <= 16'h0000;
            14'h3bde: oData <= 16'h0000;
            14'h3bdf: oData <= 16'h0000;
            14'h3be0: oData <= 16'h0000;
            14'h3be1: oData <= 16'h0000;
            14'h3be2: oData <= 16'h0000;
            14'h3be3: oData <= 16'h0000;
            14'h3be4: oData <= 16'h0000;
            14'h3be5: oData <= 16'h0000;
            14'h3be6: oData <= 16'h0000;
            14'h3be7: oData <= 16'h0000;
            14'h3be8: oData <= 16'h0000;
            14'h3be9: oData <= 16'h0000;
            14'h3bea: oData <= 16'h0000;
            14'h3beb: oData <= 16'h0000;
            14'h3bec: oData <= 16'h0000;
            14'h3bed: oData <= 16'h0000;
            14'h3bee: oData <= 16'h0000;
            14'h3bef: oData <= 16'h0000;
            14'h3bf0: oData <= 16'h0000;
            14'h3bf1: oData <= 16'h0000;
            14'h3bf2: oData <= 16'h0000;
            14'h3bf3: oData <= 16'h0000;
            14'h3bf4: oData <= 16'h0000;
            14'h3bf5: oData <= 16'h0000;
            14'h3bf6: oData <= 16'h0000;
            14'h3bf7: oData <= 16'h0000;
            14'h3bf8: oData <= 16'h0000;
            14'h3bf9: oData <= 16'h0000;
            14'h3bfa: oData <= 16'h0000;
            14'h3bfb: oData <= 16'h0000;
            14'h3bfc: oData <= 16'h0000;
            14'h3bfd: oData <= 16'h0000;
            14'h3bfe: oData <= 16'h0000;
            14'h3bff: oData <= 16'h0000;
            14'h3c00: oData <= 16'h0000;
            14'h3c01: oData <= 16'h0000;
            14'h3c02: oData <= 16'h0000;
            14'h3c03: oData <= 16'h0000;
            14'h3c04: oData <= 16'h0000;
            14'h3c05: oData <= 16'h0000;
            14'h3c06: oData <= 16'h0000;
            14'h3c07: oData <= 16'h0000;
            14'h3c08: oData <= 16'h0000;
            14'h3c09: oData <= 16'h0000;
            14'h3c0a: oData <= 16'h0000;
            14'h3c0b: oData <= 16'h0000;
            14'h3c0c: oData <= 16'h0000;
            14'h3c0d: oData <= 16'h0000;
            14'h3c0e: oData <= 16'h0000;
            14'h3c0f: oData <= 16'h0000;
            14'h3c10: oData <= 16'h0000;
            14'h3c11: oData <= 16'h0000;
            14'h3c12: oData <= 16'h0000;
            14'h3c13: oData <= 16'h0000;
            14'h3c14: oData <= 16'h0000;
            14'h3c15: oData <= 16'h0000;
            14'h3c16: oData <= 16'h0000;
            14'h3c17: oData <= 16'h0000;
            14'h3c18: oData <= 16'h0000;
            14'h3c19: oData <= 16'h0000;
            14'h3c1a: oData <= 16'h0000;
            14'h3c1b: oData <= 16'h0000;
            14'h3c1c: oData <= 16'h0000;
            14'h3c1d: oData <= 16'h0000;
            14'h3c1e: oData <= 16'h0000;
            14'h3c1f: oData <= 16'h0000;
            14'h3c20: oData <= 16'h0000;
            14'h3c21: oData <= 16'h0000;
            14'h3c22: oData <= 16'h0000;
            14'h3c23: oData <= 16'h0000;
            14'h3c24: oData <= 16'h0000;
            14'h3c25: oData <= 16'h0000;
            14'h3c26: oData <= 16'h0000;
            14'h3c27: oData <= 16'h0000;
            14'h3c28: oData <= 16'h0000;
            14'h3c29: oData <= 16'h0000;
            14'h3c2a: oData <= 16'h0000;
            14'h3c2b: oData <= 16'h0000;
            14'h3c2c: oData <= 16'h0000;
            14'h3c2d: oData <= 16'h0000;
            14'h3c2e: oData <= 16'h0000;
            14'h3c2f: oData <= 16'h0000;
            14'h3c30: oData <= 16'h0000;
            14'h3c31: oData <= 16'h0000;
            14'h3c32: oData <= 16'h0000;
            14'h3c33: oData <= 16'h0000;
            14'h3c34: oData <= 16'h0000;
            14'h3c35: oData <= 16'h0000;
            14'h3c36: oData <= 16'h0000;
            14'h3c37: oData <= 16'h0000;
            14'h3c38: oData <= 16'h0000;
            14'h3c39: oData <= 16'h0000;
            14'h3c3a: oData <= 16'h0000;
            14'h3c3b: oData <= 16'h0000;
            14'h3c3c: oData <= 16'h0000;
            14'h3c3d: oData <= 16'h0000;
            14'h3c3e: oData <= 16'h0000;
            14'h3c3f: oData <= 16'h0000;
            14'h3c40: oData <= 16'h0000;
            14'h3c41: oData <= 16'h0000;
            14'h3c42: oData <= 16'h0000;
            14'h3c43: oData <= 16'h0000;
            14'h3c44: oData <= 16'h0000;
            14'h3c45: oData <= 16'h0000;
            14'h3c46: oData <= 16'h0000;
            14'h3c47: oData <= 16'h0000;
            14'h3c48: oData <= 16'h0000;
            14'h3c49: oData <= 16'h0000;
            14'h3c4a: oData <= 16'h0000;
            14'h3c4b: oData <= 16'h0000;
            14'h3c4c: oData <= 16'h0000;
            14'h3c4d: oData <= 16'h0000;
            14'h3c4e: oData <= 16'h0000;
            14'h3c4f: oData <= 16'h0000;
            14'h3c50: oData <= 16'h0000;
            14'h3c51: oData <= 16'h0000;
            14'h3c52: oData <= 16'h0000;
            14'h3c53: oData <= 16'h0000;
            14'h3c54: oData <= 16'h0000;
            14'h3c55: oData <= 16'h0000;
            14'h3c56: oData <= 16'h0000;
            14'h3c57: oData <= 16'h0000;
            14'h3c58: oData <= 16'h0000;
            14'h3c59: oData <= 16'h0000;
            14'h3c5a: oData <= 16'h0000;
            14'h3c5b: oData <= 16'h0000;
            14'h3c5c: oData <= 16'h0000;
            14'h3c5d: oData <= 16'h0000;
            14'h3c5e: oData <= 16'h0000;
            14'h3c5f: oData <= 16'h0000;
            14'h3c60: oData <= 16'h0000;
            14'h3c61: oData <= 16'h0000;
            14'h3c62: oData <= 16'h0000;
            14'h3c63: oData <= 16'h0000;
            14'h3c64: oData <= 16'h0000;
            14'h3c65: oData <= 16'h0000;
            14'h3c66: oData <= 16'h0000;
            14'h3c67: oData <= 16'h0000;
            14'h3c68: oData <= 16'h0000;
            14'h3c69: oData <= 16'h0000;
            14'h3c6a: oData <= 16'h0000;
            14'h3c6b: oData <= 16'h0000;
            14'h3c6c: oData <= 16'h0000;
            14'h3c6d: oData <= 16'h0000;
            14'h3c6e: oData <= 16'h0000;
            14'h3c6f: oData <= 16'h0000;
            14'h3c70: oData <= 16'h0000;
            14'h3c71: oData <= 16'h0000;
            14'h3c72: oData <= 16'h0000;
            14'h3c73: oData <= 16'h0000;
            14'h3c74: oData <= 16'h0000;
            14'h3c75: oData <= 16'h0000;
            14'h3c76: oData <= 16'h0000;
            14'h3c77: oData <= 16'h0000;
            14'h3c78: oData <= 16'h0000;
            14'h3c79: oData <= 16'h0000;
            14'h3c7a: oData <= 16'h0000;
            14'h3c7b: oData <= 16'h0000;
            14'h3c7c: oData <= 16'h0000;
            14'h3c7d: oData <= 16'h0000;
            14'h3c7e: oData <= 16'h0000;
            14'h3c7f: oData <= 16'h0000;
            14'h3c80: oData <= 16'h0000;
            14'h3c81: oData <= 16'h0000;
            14'h3c82: oData <= 16'h0000;
            14'h3c83: oData <= 16'h0000;
            14'h3c84: oData <= 16'h0000;
            14'h3c85: oData <= 16'h0000;
            14'h3c86: oData <= 16'h0000;
            14'h3c87: oData <= 16'h0000;
            14'h3c88: oData <= 16'h0000;
            14'h3c89: oData <= 16'h0000;
            14'h3c8a: oData <= 16'h0000;
            14'h3c8b: oData <= 16'h0000;
            14'h3c8c: oData <= 16'h0000;
            14'h3c8d: oData <= 16'h0000;
            14'h3c8e: oData <= 16'h0000;
            14'h3c8f: oData <= 16'h0000;
            14'h3c90: oData <= 16'h0000;
            14'h3c91: oData <= 16'h0000;
            14'h3c92: oData <= 16'h0000;
            14'h3c93: oData <= 16'h0000;
            14'h3c94: oData <= 16'h0000;
            14'h3c95: oData <= 16'h0000;
            14'h3c96: oData <= 16'h0000;
            14'h3c97: oData <= 16'h0000;
            14'h3c98: oData <= 16'h0000;
            14'h3c99: oData <= 16'h0000;
            14'h3c9a: oData <= 16'h0000;
            14'h3c9b: oData <= 16'h0000;
            14'h3c9c: oData <= 16'h0000;
            14'h3c9d: oData <= 16'h0000;
            14'h3c9e: oData <= 16'h0000;
            14'h3c9f: oData <= 16'h0000;
            14'h3ca0: oData <= 16'h0000;
            14'h3ca1: oData <= 16'h0000;
            14'h3ca2: oData <= 16'h0000;
            14'h3ca3: oData <= 16'h0000;
            14'h3ca4: oData <= 16'h0000;
            14'h3ca5: oData <= 16'h0000;
            14'h3ca6: oData <= 16'h0000;
            14'h3ca7: oData <= 16'h0000;
            14'h3ca8: oData <= 16'h0000;
            14'h3ca9: oData <= 16'h0000;
            14'h3caa: oData <= 16'h0000;
            14'h3cab: oData <= 16'h0000;
            14'h3cac: oData <= 16'h0000;
            14'h3cad: oData <= 16'h0000;
            14'h3cae: oData <= 16'h0000;
            14'h3caf: oData <= 16'h0000;
            14'h3cb0: oData <= 16'h0000;
            14'h3cb1: oData <= 16'h0000;
            14'h3cb2: oData <= 16'h0000;
            14'h3cb3: oData <= 16'h0000;
            14'h3cb4: oData <= 16'h0000;
            14'h3cb5: oData <= 16'h0000;
            14'h3cb6: oData <= 16'h0000;
            14'h3cb7: oData <= 16'h0000;
            14'h3cb8: oData <= 16'h0000;
            14'h3cb9: oData <= 16'h0000;
            14'h3cba: oData <= 16'h0000;
            14'h3cbb: oData <= 16'h0000;
            14'h3cbc: oData <= 16'h0000;
            14'h3cbd: oData <= 16'h0000;
            14'h3cbe: oData <= 16'h0000;
            14'h3cbf: oData <= 16'h0000;
            14'h3cc0: oData <= 16'h0000;
            14'h3cc1: oData <= 16'h0000;
            14'h3cc2: oData <= 16'h0000;
            14'h3cc3: oData <= 16'h0000;
            14'h3cc4: oData <= 16'h0000;
            14'h3cc5: oData <= 16'h0000;
            14'h3cc6: oData <= 16'h0000;
            14'h3cc7: oData <= 16'h0000;
            14'h3cc8: oData <= 16'h0000;
            14'h3cc9: oData <= 16'h0000;
            14'h3cca: oData <= 16'h0000;
            14'h3ccb: oData <= 16'h0000;
            14'h3ccc: oData <= 16'h0000;
            14'h3ccd: oData <= 16'h0000;
            14'h3cce: oData <= 16'h0000;
            14'h3ccf: oData <= 16'h0000;
            14'h3cd0: oData <= 16'h0000;
            14'h3cd1: oData <= 16'h0000;
            14'h3cd2: oData <= 16'h0000;
            14'h3cd3: oData <= 16'h0000;
            14'h3cd4: oData <= 16'h0000;
            14'h3cd5: oData <= 16'h0000;
            14'h3cd6: oData <= 16'h0000;
            14'h3cd7: oData <= 16'h0000;
            14'h3cd8: oData <= 16'h0000;
            14'h3cd9: oData <= 16'h0000;
            14'h3cda: oData <= 16'h0000;
            14'h3cdb: oData <= 16'h0000;
            14'h3cdc: oData <= 16'h0000;
            14'h3cdd: oData <= 16'h0000;
            14'h3cde: oData <= 16'h0000;
            14'h3cdf: oData <= 16'h0000;
            14'h3ce0: oData <= 16'h0000;
            14'h3ce1: oData <= 16'h0000;
            14'h3ce2: oData <= 16'h0000;
            14'h3ce3: oData <= 16'h0000;
            14'h3ce4: oData <= 16'h0000;
            14'h3ce5: oData <= 16'h0000;
            14'h3ce6: oData <= 16'h0000;
            14'h3ce7: oData <= 16'h0000;
            14'h3ce8: oData <= 16'h0000;
            14'h3ce9: oData <= 16'h0000;
            14'h3cea: oData <= 16'h0000;
            14'h3ceb: oData <= 16'h0000;
            14'h3cec: oData <= 16'h0000;
            14'h3ced: oData <= 16'h0000;
            14'h3cee: oData <= 16'h0000;
            14'h3cef: oData <= 16'h0000;
            14'h3cf0: oData <= 16'h0000;
            14'h3cf1: oData <= 16'h0000;
            14'h3cf2: oData <= 16'h0000;
            14'h3cf3: oData <= 16'h0000;
            14'h3cf4: oData <= 16'h0000;
            14'h3cf5: oData <= 16'h0000;
            14'h3cf6: oData <= 16'h0000;
            14'h3cf7: oData <= 16'h0000;
            14'h3cf8: oData <= 16'h0000;
            14'h3cf9: oData <= 16'h0000;
            14'h3cfa: oData <= 16'h0000;
            14'h3cfb: oData <= 16'h0000;
            14'h3cfc: oData <= 16'h0000;
            14'h3cfd: oData <= 16'h0000;
            14'h3cfe: oData <= 16'h0000;
            14'h3cff: oData <= 16'h0000;
            14'h3d00: oData <= 16'h0000;
            14'h3d01: oData <= 16'h0000;
            14'h3d02: oData <= 16'h0000;
            14'h3d03: oData <= 16'h0000;
            14'h3d04: oData <= 16'h0000;
            14'h3d05: oData <= 16'h0000;
            14'h3d06: oData <= 16'h0000;
            14'h3d07: oData <= 16'h0000;
            14'h3d08: oData <= 16'h0000;
            14'h3d09: oData <= 16'h0000;
            14'h3d0a: oData <= 16'h0000;
            14'h3d0b: oData <= 16'h0000;
            14'h3d0c: oData <= 16'h0000;
            14'h3d0d: oData <= 16'h0000;
            14'h3d0e: oData <= 16'h0000;
            14'h3d0f: oData <= 16'h0000;
            14'h3d10: oData <= 16'h0000;
            14'h3d11: oData <= 16'h0000;
            14'h3d12: oData <= 16'h0000;
            14'h3d13: oData <= 16'h0000;
            14'h3d14: oData <= 16'h0000;
            14'h3d15: oData <= 16'h0000;
            14'h3d16: oData <= 16'h0000;
            14'h3d17: oData <= 16'h0000;
            14'h3d18: oData <= 16'h0000;
            14'h3d19: oData <= 16'h0000;
            14'h3d1a: oData <= 16'h0000;
            14'h3d1b: oData <= 16'h0000;
            14'h3d1c: oData <= 16'h0000;
            14'h3d1d: oData <= 16'h0000;
            14'h3d1e: oData <= 16'h0000;
            14'h3d1f: oData <= 16'h0000;
            14'h3d20: oData <= 16'h0000;
            14'h3d21: oData <= 16'h0000;
            14'h3d22: oData <= 16'h0000;
            14'h3d23: oData <= 16'h0000;
            14'h3d24: oData <= 16'h0000;
            14'h3d25: oData <= 16'h0000;
            14'h3d26: oData <= 16'h0000;
            14'h3d27: oData <= 16'h0000;
            14'h3d28: oData <= 16'h0000;
            14'h3d29: oData <= 16'h0000;
            14'h3d2a: oData <= 16'h0000;
            14'h3d2b: oData <= 16'h0000;
            14'h3d2c: oData <= 16'h0000;
            14'h3d2d: oData <= 16'h0000;
            14'h3d2e: oData <= 16'h0000;
            14'h3d2f: oData <= 16'h0000;
            14'h3d30: oData <= 16'h0000;
            14'h3d31: oData <= 16'h0000;
            14'h3d32: oData <= 16'h0000;
            14'h3d33: oData <= 16'h0000;
            14'h3d34: oData <= 16'h0000;
            14'h3d35: oData <= 16'h0000;
            14'h3d36: oData <= 16'h0000;
            14'h3d37: oData <= 16'h0000;
            14'h3d38: oData <= 16'h0000;
            14'h3d39: oData <= 16'h0000;
            14'h3d3a: oData <= 16'h0000;
            14'h3d3b: oData <= 16'h0000;
            14'h3d3c: oData <= 16'h0000;
            14'h3d3d: oData <= 16'h0000;
            14'h3d3e: oData <= 16'h0000;
            14'h3d3f: oData <= 16'h0000;
            14'h3d40: oData <= 16'h0000;
            14'h3d41: oData <= 16'h0000;
            14'h3d42: oData <= 16'h0000;
            14'h3d43: oData <= 16'h0000;
            14'h3d44: oData <= 16'h0000;
            14'h3d45: oData <= 16'h0000;
            14'h3d46: oData <= 16'h0000;
            14'h3d47: oData <= 16'h0000;
            14'h3d48: oData <= 16'h0000;
            14'h3d49: oData <= 16'h0000;
            14'h3d4a: oData <= 16'h0000;
            14'h3d4b: oData <= 16'h0000;
            14'h3d4c: oData <= 16'h0000;
            14'h3d4d: oData <= 16'h0000;
            14'h3d4e: oData <= 16'h0000;
            14'h3d4f: oData <= 16'h0000;
            14'h3d50: oData <= 16'h0000;
            14'h3d51: oData <= 16'h0000;
            14'h3d52: oData <= 16'h0000;
            14'h3d53: oData <= 16'h0000;
            14'h3d54: oData <= 16'h0000;
            14'h3d55: oData <= 16'h0000;
            14'h3d56: oData <= 16'h0000;
            14'h3d57: oData <= 16'h0000;
            14'h3d58: oData <= 16'h0000;
            14'h3d59: oData <= 16'h0000;
            14'h3d5a: oData <= 16'h0000;
            14'h3d5b: oData <= 16'h0000;
            14'h3d5c: oData <= 16'h0000;
            14'h3d5d: oData <= 16'h0000;
            14'h3d5e: oData <= 16'h0000;
            14'h3d5f: oData <= 16'h0000;
            14'h3d60: oData <= 16'h0000;
            14'h3d61: oData <= 16'h0000;
            14'h3d62: oData <= 16'h0000;
            14'h3d63: oData <= 16'h0000;
            14'h3d64: oData <= 16'h0000;
            14'h3d65: oData <= 16'h0000;
            14'h3d66: oData <= 16'h0000;
            14'h3d67: oData <= 16'h0000;
            14'h3d68: oData <= 16'h0000;
            14'h3d69: oData <= 16'h0000;
            14'h3d6a: oData <= 16'h0000;
            14'h3d6b: oData <= 16'h0000;
            14'h3d6c: oData <= 16'h0000;
            14'h3d6d: oData <= 16'h0000;
            14'h3d6e: oData <= 16'h0000;
            14'h3d6f: oData <= 16'h0000;
            14'h3d70: oData <= 16'h0000;
            14'h3d71: oData <= 16'h0000;
            14'h3d72: oData <= 16'h0000;
            14'h3d73: oData <= 16'h0000;
            14'h3d74: oData <= 16'h0000;
            14'h3d75: oData <= 16'h0000;
            14'h3d76: oData <= 16'h0000;
            14'h3d77: oData <= 16'h0000;
            14'h3d78: oData <= 16'h0000;
            14'h3d79: oData <= 16'h0000;
            14'h3d7a: oData <= 16'h0000;
            14'h3d7b: oData <= 16'h0000;
            14'h3d7c: oData <= 16'h0000;
            14'h3d7d: oData <= 16'h0000;
            14'h3d7e: oData <= 16'h0000;
            14'h3d7f: oData <= 16'h0000;
            14'h3d80: oData <= 16'h0000;
            14'h3d81: oData <= 16'h0000;
            14'h3d82: oData <= 16'h0000;
            14'h3d83: oData <= 16'h0000;
            14'h3d84: oData <= 16'h0000;
            14'h3d85: oData <= 16'h0000;
            14'h3d86: oData <= 16'h0000;
            14'h3d87: oData <= 16'h0000;
            14'h3d88: oData <= 16'h0000;
            14'h3d89: oData <= 16'h0000;
            14'h3d8a: oData <= 16'h0000;
            14'h3d8b: oData <= 16'h0000;
            14'h3d8c: oData <= 16'h0000;
            14'h3d8d: oData <= 16'h0000;
            14'h3d8e: oData <= 16'h0000;
            14'h3d8f: oData <= 16'h0000;
            14'h3d90: oData <= 16'h0000;
            14'h3d91: oData <= 16'h0000;
            14'h3d92: oData <= 16'h0000;
            14'h3d93: oData <= 16'h0000;
            14'h3d94: oData <= 16'h0000;
            14'h3d95: oData <= 16'h0000;
            14'h3d96: oData <= 16'h0000;
            14'h3d97: oData <= 16'h0000;
            14'h3d98: oData <= 16'h0000;
            14'h3d99: oData <= 16'h0000;
            14'h3d9a: oData <= 16'h0000;
            14'h3d9b: oData <= 16'h0000;
            14'h3d9c: oData <= 16'h0000;
            14'h3d9d: oData <= 16'h0000;
            14'h3d9e: oData <= 16'h0000;
            14'h3d9f: oData <= 16'h0000;
            14'h3da0: oData <= 16'h0000;
            14'h3da1: oData <= 16'h0000;
            14'h3da2: oData <= 16'h0000;
            14'h3da3: oData <= 16'h0000;
            14'h3da4: oData <= 16'h0000;
            14'h3da5: oData <= 16'h0000;
            14'h3da6: oData <= 16'h0000;
            14'h3da7: oData <= 16'h0000;
            14'h3da8: oData <= 16'h0000;
            14'h3da9: oData <= 16'h0000;
            14'h3daa: oData <= 16'h0000;
            14'h3dab: oData <= 16'h0000;
            14'h3dac: oData <= 16'h0000;
            14'h3dad: oData <= 16'h0000;
            14'h3dae: oData <= 16'h0000;
            14'h3daf: oData <= 16'h0000;
            14'h3db0: oData <= 16'h0000;
            14'h3db1: oData <= 16'h0000;
            14'h3db2: oData <= 16'h0000;
            14'h3db3: oData <= 16'h0000;
            14'h3db4: oData <= 16'h0000;
            14'h3db5: oData <= 16'h0000;
            14'h3db6: oData <= 16'h0000;
            14'h3db7: oData <= 16'h0000;
            14'h3db8: oData <= 16'h0000;
            14'h3db9: oData <= 16'h0000;
            14'h3dba: oData <= 16'h0000;
            14'h3dbb: oData <= 16'h0000;
            14'h3dbc: oData <= 16'h0000;
            14'h3dbd: oData <= 16'h0000;
            14'h3dbe: oData <= 16'h0000;
            14'h3dbf: oData <= 16'h0000;
            14'h3dc0: oData <= 16'h0000;
            14'h3dc1: oData <= 16'h0000;
            14'h3dc2: oData <= 16'h0000;
            14'h3dc3: oData <= 16'h0000;
            14'h3dc4: oData <= 16'h0000;
            14'h3dc5: oData <= 16'h0000;
            14'h3dc6: oData <= 16'h0000;
            14'h3dc7: oData <= 16'h0000;
            14'h3dc8: oData <= 16'h0000;
            14'h3dc9: oData <= 16'h0000;
            14'h3dca: oData <= 16'h0000;
            14'h3dcb: oData <= 16'h0000;
            14'h3dcc: oData <= 16'h0000;
            14'h3dcd: oData <= 16'h0000;
            14'h3dce: oData <= 16'h0000;
            14'h3dcf: oData <= 16'h0000;
            14'h3dd0: oData <= 16'h0000;
            14'h3dd1: oData <= 16'h0000;
            14'h3dd2: oData <= 16'h0000;
            14'h3dd3: oData <= 16'h0000;
            14'h3dd4: oData <= 16'h0000;
            14'h3dd5: oData <= 16'h0000;
            14'h3dd6: oData <= 16'h0000;
            14'h3dd7: oData <= 16'h0000;
            14'h3dd8: oData <= 16'h0000;
            14'h3dd9: oData <= 16'h0000;
            14'h3dda: oData <= 16'h0000;
            14'h3ddb: oData <= 16'h0000;
            14'h3ddc: oData <= 16'h0000;
            14'h3ddd: oData <= 16'h0000;
            14'h3dde: oData <= 16'h0000;
            14'h3ddf: oData <= 16'h0000;
            14'h3de0: oData <= 16'h0000;
            14'h3de1: oData <= 16'h0000;
            14'h3de2: oData <= 16'h0000;
            14'h3de3: oData <= 16'h0000;
            14'h3de4: oData <= 16'h0000;
            14'h3de5: oData <= 16'h0000;
            14'h3de6: oData <= 16'h0000;
            14'h3de7: oData <= 16'h0000;
            14'h3de8: oData <= 16'h0000;
            14'h3de9: oData <= 16'h0000;
            14'h3dea: oData <= 16'h0000;
            14'h3deb: oData <= 16'h0000;
            14'h3dec: oData <= 16'h0000;
            14'h3ded: oData <= 16'h0000;
            14'h3dee: oData <= 16'h0000;
            14'h3def: oData <= 16'h0000;
            14'h3df0: oData <= 16'h0000;
            14'h3df1: oData <= 16'h0000;
            14'h3df2: oData <= 16'h0000;
            14'h3df3: oData <= 16'h0000;
            14'h3df4: oData <= 16'h0000;
            14'h3df5: oData <= 16'h0000;
            14'h3df6: oData <= 16'h0000;
            14'h3df7: oData <= 16'h0000;
            14'h3df8: oData <= 16'h0000;
            14'h3df9: oData <= 16'h0000;
            14'h3dfa: oData <= 16'h0000;
            14'h3dfb: oData <= 16'h0000;
            14'h3dfc: oData <= 16'h0000;
            14'h3dfd: oData <= 16'h0000;
            14'h3dfe: oData <= 16'h0000;
            14'h3dff: oData <= 16'h0000;
            14'h3e00: oData <= 16'h0000;
            14'h3e01: oData <= 16'h0000;
            14'h3e02: oData <= 16'h0000;
            14'h3e03: oData <= 16'h0000;
            14'h3e04: oData <= 16'h0000;
            14'h3e05: oData <= 16'h0000;
            14'h3e06: oData <= 16'h0000;
            14'h3e07: oData <= 16'h0000;
            14'h3e08: oData <= 16'h0000;
            14'h3e09: oData <= 16'h0000;
            14'h3e0a: oData <= 16'h0000;
            14'h3e0b: oData <= 16'h0000;
            14'h3e0c: oData <= 16'h0000;
            14'h3e0d: oData <= 16'h0000;
            14'h3e0e: oData <= 16'h0000;
            14'h3e0f: oData <= 16'h0000;
            14'h3e10: oData <= 16'h0000;
            14'h3e11: oData <= 16'h0000;
            14'h3e12: oData <= 16'h0000;
            14'h3e13: oData <= 16'h0000;
            14'h3e14: oData <= 16'h0000;
            14'h3e15: oData <= 16'h0000;
            14'h3e16: oData <= 16'h0000;
            14'h3e17: oData <= 16'h0000;
            14'h3e18: oData <= 16'h0000;
            14'h3e19: oData <= 16'h0000;
            14'h3e1a: oData <= 16'h0000;
            14'h3e1b: oData <= 16'h0000;
            14'h3e1c: oData <= 16'h0000;
            14'h3e1d: oData <= 16'h0000;
            14'h3e1e: oData <= 16'h0000;
            14'h3e1f: oData <= 16'h0000;
            14'h3e20: oData <= 16'h0000;
            14'h3e21: oData <= 16'h0000;
            14'h3e22: oData <= 16'h0000;
            14'h3e23: oData <= 16'h0000;
            14'h3e24: oData <= 16'h0000;
            14'h3e25: oData <= 16'h0000;
            14'h3e26: oData <= 16'h0000;
            14'h3e27: oData <= 16'h0000;
            14'h3e28: oData <= 16'h0000;
            14'h3e29: oData <= 16'h0000;
            14'h3e2a: oData <= 16'h0000;
            14'h3e2b: oData <= 16'h0000;
            14'h3e2c: oData <= 16'h0000;
            14'h3e2d: oData <= 16'h0000;
            14'h3e2e: oData <= 16'h0000;
            14'h3e2f: oData <= 16'h0000;
            14'h3e30: oData <= 16'h0000;
            14'h3e31: oData <= 16'h0000;
            14'h3e32: oData <= 16'h0000;
            14'h3e33: oData <= 16'h0000;
            14'h3e34: oData <= 16'h0000;
            14'h3e35: oData <= 16'h0000;
            14'h3e36: oData <= 16'h0000;
            14'h3e37: oData <= 16'h0000;
            14'h3e38: oData <= 16'h0000;
            14'h3e39: oData <= 16'h0000;
            14'h3e3a: oData <= 16'h0000;
            14'h3e3b: oData <= 16'h0000;
            14'h3e3c: oData <= 16'h0000;
            14'h3e3d: oData <= 16'h0000;
            14'h3e3e: oData <= 16'h0000;
            14'h3e3f: oData <= 16'h0000;
            14'h3e40: oData <= 16'h0000;
            14'h3e41: oData <= 16'h0000;
            14'h3e42: oData <= 16'h0000;
            14'h3e43: oData <= 16'h0000;
            14'h3e44: oData <= 16'h0000;
            14'h3e45: oData <= 16'h0000;
            14'h3e46: oData <= 16'h0000;
            14'h3e47: oData <= 16'h0000;
            14'h3e48: oData <= 16'h0000;
            14'h3e49: oData <= 16'h0000;
            14'h3e4a: oData <= 16'h0000;
            14'h3e4b: oData <= 16'h0000;
            14'h3e4c: oData <= 16'h0000;
            14'h3e4d: oData <= 16'h0000;
            14'h3e4e: oData <= 16'h0000;
            14'h3e4f: oData <= 16'h0000;
            14'h3e50: oData <= 16'h0000;
            14'h3e51: oData <= 16'h0000;
            14'h3e52: oData <= 16'h0000;
            14'h3e53: oData <= 16'h0000;
            14'h3e54: oData <= 16'h0000;
            14'h3e55: oData <= 16'h0000;
            14'h3e56: oData <= 16'h0000;
            14'h3e57: oData <= 16'h0000;
            14'h3e58: oData <= 16'h0000;
            14'h3e59: oData <= 16'h0000;
            14'h3e5a: oData <= 16'h0000;
            14'h3e5b: oData <= 16'h0000;
            14'h3e5c: oData <= 16'h0000;
            14'h3e5d: oData <= 16'h0000;
            14'h3e5e: oData <= 16'h0000;
            14'h3e5f: oData <= 16'h0000;
            14'h3e60: oData <= 16'h0000;
            14'h3e61: oData <= 16'h0000;
            14'h3e62: oData <= 16'h0000;
            14'h3e63: oData <= 16'h0000;
            14'h3e64: oData <= 16'h0000;
            14'h3e65: oData <= 16'h0000;
            14'h3e66: oData <= 16'h0000;
            14'h3e67: oData <= 16'h0000;
            14'h3e68: oData <= 16'h0000;
            14'h3e69: oData <= 16'h0000;
            14'h3e6a: oData <= 16'h0000;
            14'h3e6b: oData <= 16'h0000;
            14'h3e6c: oData <= 16'h0000;
            14'h3e6d: oData <= 16'h0000;
            14'h3e6e: oData <= 16'h0000;
            14'h3e6f: oData <= 16'h0000;
            14'h3e70: oData <= 16'h0000;
            14'h3e71: oData <= 16'h0000;
            14'h3e72: oData <= 16'h0000;
            14'h3e73: oData <= 16'h0000;
            14'h3e74: oData <= 16'h0000;
            14'h3e75: oData <= 16'h0000;
            14'h3e76: oData <= 16'h0000;
            14'h3e77: oData <= 16'h0000;
            14'h3e78: oData <= 16'h0000;
            14'h3e79: oData <= 16'h0000;
            14'h3e7a: oData <= 16'h0000;
            14'h3e7b: oData <= 16'h0000;
            14'h3e7c: oData <= 16'h0000;
            14'h3e7d: oData <= 16'h0000;
            14'h3e7e: oData <= 16'h0000;
            14'h3e7f: oData <= 16'h0000;
            14'h3e80: oData <= 16'h0000;
            14'h3e81: oData <= 16'h0000;
            14'h3e82: oData <= 16'h0000;
            14'h3e83: oData <= 16'h0000;
            14'h3e84: oData <= 16'h0000;
            14'h3e85: oData <= 16'h0000;
            14'h3e86: oData <= 16'h0000;
            14'h3e87: oData <= 16'h0000;
            14'h3e88: oData <= 16'h0000;
            14'h3e89: oData <= 16'h0000;
            14'h3e8a: oData <= 16'h0000;
            14'h3e8b: oData <= 16'h0000;
            14'h3e8c: oData <= 16'h0000;
            14'h3e8d: oData <= 16'h0000;
            14'h3e8e: oData <= 16'h0000;
            14'h3e8f: oData <= 16'h0000;
            14'h3e90: oData <= 16'h0000;
            14'h3e91: oData <= 16'h0000;
            14'h3e92: oData <= 16'h0000;
            14'h3e93: oData <= 16'h0000;
            14'h3e94: oData <= 16'h0000;
            14'h3e95: oData <= 16'h0000;
            14'h3e96: oData <= 16'h0000;
            14'h3e97: oData <= 16'h0000;
            14'h3e98: oData <= 16'h0000;
            14'h3e99: oData <= 16'h0000;
            14'h3e9a: oData <= 16'h0000;
            14'h3e9b: oData <= 16'h0000;
            14'h3e9c: oData <= 16'h0000;
            14'h3e9d: oData <= 16'h0000;
            14'h3e9e: oData <= 16'h0000;
            14'h3e9f: oData <= 16'h0000;
            14'h3ea0: oData <= 16'h0000;
            14'h3ea1: oData <= 16'h0000;
            14'h3ea2: oData <= 16'h0000;
            14'h3ea3: oData <= 16'h0000;
            14'h3ea4: oData <= 16'h0000;
            14'h3ea5: oData <= 16'h0000;
            14'h3ea6: oData <= 16'h0000;
            14'h3ea7: oData <= 16'h0000;
            14'h3ea8: oData <= 16'h0000;
            14'h3ea9: oData <= 16'h0000;
            14'h3eaa: oData <= 16'h0000;
            14'h3eab: oData <= 16'h0000;
            14'h3eac: oData <= 16'h0000;
            14'h3ead: oData <= 16'h0000;
            14'h3eae: oData <= 16'h0000;
            14'h3eaf: oData <= 16'h0000;
            14'h3eb0: oData <= 16'h0000;
            14'h3eb1: oData <= 16'h0000;
            14'h3eb2: oData <= 16'h0000;
            14'h3eb3: oData <= 16'h0000;
            14'h3eb4: oData <= 16'h0000;
            14'h3eb5: oData <= 16'h0000;
            14'h3eb6: oData <= 16'h0000;
            14'h3eb7: oData <= 16'h0000;
            14'h3eb8: oData <= 16'h0000;
            14'h3eb9: oData <= 16'h0000;
            14'h3eba: oData <= 16'h0000;
            14'h3ebb: oData <= 16'h0000;
            14'h3ebc: oData <= 16'h0000;
            14'h3ebd: oData <= 16'h0000;
            14'h3ebe: oData <= 16'h0000;
            14'h3ebf: oData <= 16'h0000;
            14'h3ec0: oData <= 16'h0000;
            14'h3ec1: oData <= 16'h0000;
            14'h3ec2: oData <= 16'h0000;
            14'h3ec3: oData <= 16'h0000;
            14'h3ec4: oData <= 16'h0000;
            14'h3ec5: oData <= 16'h0000;
            14'h3ec6: oData <= 16'h0000;
            14'h3ec7: oData <= 16'h0000;
            14'h3ec8: oData <= 16'h0000;
            14'h3ec9: oData <= 16'h0000;
            14'h3eca: oData <= 16'h0000;
            14'h3ecb: oData <= 16'h0000;
            14'h3ecc: oData <= 16'h0000;
            14'h3ecd: oData <= 16'h0000;
            14'h3ece: oData <= 16'h0000;
            14'h3ecf: oData <= 16'h0000;
            14'h3ed0: oData <= 16'h0000;
            14'h3ed1: oData <= 16'h0000;
            14'h3ed2: oData <= 16'h0000;
            14'h3ed3: oData <= 16'h0000;
            14'h3ed4: oData <= 16'h0000;
            14'h3ed5: oData <= 16'h0000;
            14'h3ed6: oData <= 16'h0000;
            14'h3ed7: oData <= 16'h0000;
            14'h3ed8: oData <= 16'h0000;
            14'h3ed9: oData <= 16'h0000;
            14'h3eda: oData <= 16'h0000;
            14'h3edb: oData <= 16'h0000;
            14'h3edc: oData <= 16'h0000;
            14'h3edd: oData <= 16'h0000;
            14'h3ede: oData <= 16'h0000;
            14'h3edf: oData <= 16'h0000;
            14'h3ee0: oData <= 16'h0000;
            14'h3ee1: oData <= 16'h0000;
            14'h3ee2: oData <= 16'h0000;
            14'h3ee3: oData <= 16'h0000;
            14'h3ee4: oData <= 16'h0000;
            14'h3ee5: oData <= 16'h0000;
            14'h3ee6: oData <= 16'h0000;
            14'h3ee7: oData <= 16'h0000;
            14'h3ee8: oData <= 16'h0000;
            14'h3ee9: oData <= 16'h0000;
            14'h3eea: oData <= 16'h0000;
            14'h3eeb: oData <= 16'h0000;
            14'h3eec: oData <= 16'h0000;
            14'h3eed: oData <= 16'h0000;
            14'h3eee: oData <= 16'h0000;
            14'h3eef: oData <= 16'h0000;
            14'h3ef0: oData <= 16'h0000;
            14'h3ef1: oData <= 16'h0000;
            14'h3ef2: oData <= 16'h0000;
            14'h3ef3: oData <= 16'h0000;
            14'h3ef4: oData <= 16'h0000;
            14'h3ef5: oData <= 16'h0000;
            14'h3ef6: oData <= 16'h0000;
            14'h3ef7: oData <= 16'h0000;
            14'h3ef8: oData <= 16'h0000;
            14'h3ef9: oData <= 16'h0000;
            14'h3efa: oData <= 16'h0000;
            14'h3efb: oData <= 16'h0000;
            14'h3efc: oData <= 16'h0000;
            14'h3efd: oData <= 16'h0000;
            14'h3efe: oData <= 16'h0000;
            14'h3eff: oData <= 16'h0000;
            14'h3f00: oData <= 16'h0000;
            14'h3f01: oData <= 16'h0000;
            14'h3f02: oData <= 16'h0000;
            14'h3f03: oData <= 16'h0000;
            14'h3f04: oData <= 16'h0000;
            14'h3f05: oData <= 16'h0000;
            14'h3f06: oData <= 16'h0000;
            14'h3f07: oData <= 16'h0000;
            14'h3f08: oData <= 16'h0000;
            14'h3f09: oData <= 16'h0000;
            14'h3f0a: oData <= 16'h0000;
            14'h3f0b: oData <= 16'h0000;
            14'h3f0c: oData <= 16'h0000;
            14'h3f0d: oData <= 16'h0000;
            14'h3f0e: oData <= 16'h0000;
            14'h3f0f: oData <= 16'h0000;
            14'h3f10: oData <= 16'h0000;
            14'h3f11: oData <= 16'h0000;
            14'h3f12: oData <= 16'h0000;
            14'h3f13: oData <= 16'h0000;
            14'h3f14: oData <= 16'h0000;
            14'h3f15: oData <= 16'h0000;
            14'h3f16: oData <= 16'h0000;
            14'h3f17: oData <= 16'h0000;
            14'h3f18: oData <= 16'h0000;
            14'h3f19: oData <= 16'h0000;
            14'h3f1a: oData <= 16'h0000;
            14'h3f1b: oData <= 16'h0000;
            14'h3f1c: oData <= 16'h0000;
            14'h3f1d: oData <= 16'h0000;
            14'h3f1e: oData <= 16'h0000;
            14'h3f1f: oData <= 16'h0000;
            14'h3f20: oData <= 16'h0000;
            14'h3f21: oData <= 16'h0000;
            14'h3f22: oData <= 16'h0000;
            14'h3f23: oData <= 16'h0000;
            14'h3f24: oData <= 16'h0000;
            14'h3f25: oData <= 16'h0000;
            14'h3f26: oData <= 16'h0000;
            14'h3f27: oData <= 16'h0000;
            14'h3f28: oData <= 16'h0000;
            14'h3f29: oData <= 16'h0000;
            14'h3f2a: oData <= 16'h0000;
            14'h3f2b: oData <= 16'h0000;
            14'h3f2c: oData <= 16'h0000;
            14'h3f2d: oData <= 16'h0000;
            14'h3f2e: oData <= 16'h0000;
            14'h3f2f: oData <= 16'h0000;
            14'h3f30: oData <= 16'h0000;
            14'h3f31: oData <= 16'h0000;
            14'h3f32: oData <= 16'h0000;
            14'h3f33: oData <= 16'h0000;
            14'h3f34: oData <= 16'h0000;
            14'h3f35: oData <= 16'h0000;
            14'h3f36: oData <= 16'h0000;
            14'h3f37: oData <= 16'h0000;
            14'h3f38: oData <= 16'h0000;
            14'h3f39: oData <= 16'h0000;
            14'h3f3a: oData <= 16'h0000;
            14'h3f3b: oData <= 16'h0000;
            14'h3f3c: oData <= 16'h0000;
            14'h3f3d: oData <= 16'h0000;
            14'h3f3e: oData <= 16'h0000;
            14'h3f3f: oData <= 16'h0000;
            14'h3f40: oData <= 16'h0000;
            14'h3f41: oData <= 16'h0000;
            14'h3f42: oData <= 16'h0000;
            14'h3f43: oData <= 16'h0000;
            14'h3f44: oData <= 16'h0000;
            14'h3f45: oData <= 16'h0000;
            14'h3f46: oData <= 16'h0000;
            14'h3f47: oData <= 16'h0000;
            14'h3f48: oData <= 16'h0000;
            14'h3f49: oData <= 16'h0000;
            14'h3f4a: oData <= 16'h0000;
            14'h3f4b: oData <= 16'h0000;
            14'h3f4c: oData <= 16'h0000;
            14'h3f4d: oData <= 16'h0000;
            14'h3f4e: oData <= 16'h0000;
            14'h3f4f: oData <= 16'h0000;
            14'h3f50: oData <= 16'h0000;
            14'h3f51: oData <= 16'h0000;
            14'h3f52: oData <= 16'h0000;
            14'h3f53: oData <= 16'h0000;
            14'h3f54: oData <= 16'h0000;
            14'h3f55: oData <= 16'h0000;
            14'h3f56: oData <= 16'h0000;
            14'h3f57: oData <= 16'h0000;
            14'h3f58: oData <= 16'h0000;
            14'h3f59: oData <= 16'h0000;
            14'h3f5a: oData <= 16'h0000;
            14'h3f5b: oData <= 16'h0000;
            14'h3f5c: oData <= 16'h0000;
            14'h3f5d: oData <= 16'h0000;
            14'h3f5e: oData <= 16'h0000;
            14'h3f5f: oData <= 16'h0000;
            14'h3f60: oData <= 16'h0000;
            14'h3f61: oData <= 16'h0000;
            14'h3f62: oData <= 16'h0000;
            14'h3f63: oData <= 16'h0000;
            14'h3f64: oData <= 16'h0000;
            14'h3f65: oData <= 16'h0000;
            14'h3f66: oData <= 16'h0000;
            14'h3f67: oData <= 16'h0000;
            14'h3f68: oData <= 16'h0000;
            14'h3f69: oData <= 16'h0000;
            14'h3f6a: oData <= 16'h0000;
            14'h3f6b: oData <= 16'h0000;
            14'h3f6c: oData <= 16'h0000;
            14'h3f6d: oData <= 16'h0000;
            14'h3f6e: oData <= 16'h0000;
            14'h3f6f: oData <= 16'h0000;
            14'h3f70: oData <= 16'h0000;
            14'h3f71: oData <= 16'h0000;
            14'h3f72: oData <= 16'h0000;
            14'h3f73: oData <= 16'h0000;
            14'h3f74: oData <= 16'h0000;
            14'h3f75: oData <= 16'h0000;
            14'h3f76: oData <= 16'h0000;
            14'h3f77: oData <= 16'h0000;
            14'h3f78: oData <= 16'h0000;
            14'h3f79: oData <= 16'h0000;
            14'h3f7a: oData <= 16'h0000;
            14'h3f7b: oData <= 16'h0000;
            14'h3f7c: oData <= 16'h0000;
            14'h3f7d: oData <= 16'h0000;
            14'h3f7e: oData <= 16'h0000;
            14'h3f7f: oData <= 16'h0000;
            14'h3f80: oData <= 16'h0000;
            14'h3f81: oData <= 16'h0000;
            14'h3f82: oData <= 16'h0000;
            14'h3f83: oData <= 16'h0000;
            14'h3f84: oData <= 16'h0000;
            14'h3f85: oData <= 16'h0000;
            14'h3f86: oData <= 16'h0000;
            14'h3f87: oData <= 16'h0000;
            14'h3f88: oData <= 16'h0000;
            14'h3f89: oData <= 16'h0000;
            14'h3f8a: oData <= 16'h0000;
            14'h3f8b: oData <= 16'h0000;
            14'h3f8c: oData <= 16'h0000;
            14'h3f8d: oData <= 16'h0000;
            14'h3f8e: oData <= 16'h0000;
            14'h3f8f: oData <= 16'h0000;
            14'h3f90: oData <= 16'h0000;
            14'h3f91: oData <= 16'h0000;
            14'h3f92: oData <= 16'h0000;
            14'h3f93: oData <= 16'h0000;
            14'h3f94: oData <= 16'h0000;
            14'h3f95: oData <= 16'h0000;
            14'h3f96: oData <= 16'h0000;
            14'h3f97: oData <= 16'h0000;
            14'h3f98: oData <= 16'h0000;
            14'h3f99: oData <= 16'h0000;
            14'h3f9a: oData <= 16'h0000;
            14'h3f9b: oData <= 16'h0000;
            14'h3f9c: oData <= 16'h0000;
            14'h3f9d: oData <= 16'h0000;
            14'h3f9e: oData <= 16'h0000;
            14'h3f9f: oData <= 16'h0000;
            14'h3fa0: oData <= 16'h0000;
            14'h3fa1: oData <= 16'h0000;
            14'h3fa2: oData <= 16'h0000;
            14'h3fa3: oData <= 16'h0000;
            14'h3fa4: oData <= 16'h0000;
            14'h3fa5: oData <= 16'h0000;
            14'h3fa6: oData <= 16'h0000;
            14'h3fa7: oData <= 16'h0000;
            14'h3fa8: oData <= 16'h0000;
            14'h3fa9: oData <= 16'h0000;
            14'h3faa: oData <= 16'h0000;
            14'h3fab: oData <= 16'h0000;
            14'h3fac: oData <= 16'h0000;
            14'h3fad: oData <= 16'h0000;
            14'h3fae: oData <= 16'h0000;
            14'h3faf: oData <= 16'h0000;
            14'h3fb0: oData <= 16'h0000;
            14'h3fb1: oData <= 16'h0000;
            14'h3fb2: oData <= 16'h0000;
            14'h3fb3: oData <= 16'h0000;
            14'h3fb4: oData <= 16'h0000;
            14'h3fb5: oData <= 16'h0000;
            14'h3fb6: oData <= 16'h0000;
            14'h3fb7: oData <= 16'h0000;
            14'h3fb8: oData <= 16'h0000;
            14'h3fb9: oData <= 16'h0000;
            14'h3fba: oData <= 16'h0000;
            14'h3fbb: oData <= 16'h0000;
            14'h3fbc: oData <= 16'h0000;
            14'h3fbd: oData <= 16'h0000;
            14'h3fbe: oData <= 16'h0000;
            14'h3fbf: oData <= 16'h0000;
            14'h3fc0: oData <= 16'h0000;
            14'h3fc1: oData <= 16'h0000;
            14'h3fc2: oData <= 16'h0000;
            14'h3fc3: oData <= 16'h0000;
            14'h3fc4: oData <= 16'h0000;
            14'h3fc5: oData <= 16'h0000;
            14'h3fc6: oData <= 16'h0000;
            14'h3fc7: oData <= 16'h0000;
            14'h3fc8: oData <= 16'h0000;
            14'h3fc9: oData <= 16'h0000;
            14'h3fca: oData <= 16'h0000;
            14'h3fcb: oData <= 16'h0000;
            14'h3fcc: oData <= 16'h0000;
            14'h3fcd: oData <= 16'h0000;
            14'h3fce: oData <= 16'h0000;
            14'h3fcf: oData <= 16'h0000;
            14'h3fd0: oData <= 16'h0000;
            14'h3fd1: oData <= 16'h0000;
            14'h3fd2: oData <= 16'h0000;
            14'h3fd3: oData <= 16'h0000;
            14'h3fd4: oData <= 16'h0000;
            14'h3fd5: oData <= 16'h0000;
            14'h3fd6: oData <= 16'h0000;
            14'h3fd7: oData <= 16'h0000;
            14'h3fd8: oData <= 16'h0000;
            14'h3fd9: oData <= 16'h0000;
            14'h3fda: oData <= 16'h0000;
            14'h3fdb: oData <= 16'h0000;
            14'h3fdc: oData <= 16'h0000;
            14'h3fdd: oData <= 16'h0000;
            14'h3fde: oData <= 16'h0000;
            14'h3fdf: oData <= 16'h0000;
            14'h3fe0: oData <= 16'h0000;
            14'h3fe1: oData <= 16'h0000;
            14'h3fe2: oData <= 16'h0000;
            14'h3fe3: oData <= 16'h0000;
            14'h3fe4: oData <= 16'h0000;
            14'h3fe5: oData <= 16'h0000;
            14'h3fe6: oData <= 16'h0000;
            14'h3fe7: oData <= 16'h0000;
            14'h3fe8: oData <= 16'h0000;
            14'h3fe9: oData <= 16'h0000;
            14'h3fea: oData <= 16'h0000;
            14'h3feb: oData <= 16'h0000;
            14'h3fec: oData <= 16'h0000;
            14'h3fed: oData <= 16'h0000;
            14'h3fee: oData <= 16'h0000;
            14'h3fef: oData <= 16'h0000;
            14'h3ff0: oData <= 16'h0000;
            14'h3ff1: oData <= 16'h0000;
            14'h3ff2: oData <= 16'h0000;
            14'h3ff3: oData <= 16'h0000;
            14'h3ff4: oData <= 16'h0000;
            14'h3ff5: oData <= 16'h0000;
            14'h3ff6: oData <= 16'h0000;
            14'h3ff7: oData <= 16'h0000;
            14'h3ff8: oData <= 16'h0000;
            14'h3ff9: oData <= 16'h0000;
            14'h3ffa: oData <= 16'h0000;
            14'h3ffb: oData <= 16'h0000;
            14'h3ffc: oData <= 16'h0000;
            14'h3ffd: oData <= 16'h0000;
            14'h3ffe: oData <= 16'h0000;
            14'h3fff: oData <= 16'h0000;
        endcase
    end
endmodule
