//module SEG7_LUT_8 (	oSEG0,oSEG1,oSEG2,oSEG3,oSEG4,oSEG5,oSEG6,oSEG7,iDIG );
//input	[31:0]	iDIG;
//output	[6:0]	oSEG0,oSEG1,oSEG2,oSEG3,oSEG4,oSEG5,oSEG6,oSEG7;
module SEG7_LUT_8 (	oSEG0,oSEG1,oSEG2,oSEG3,iDIG );
input	[31:0]	iDIG;
output	[6:0]	oSEG0,oSEG1,oSEG2,oSEG3;

SEG7_LUT	u0	(	oSEG0,iDIG[3:0]		);
SEG7_LUT	u1	(	oSEG1,iDIG[7:4]		);
SEG7_LUT	u2	(	oSEG2,iDIG[11:8]	);
//SEG7_LUT	u3	(	oSEG3,iDIG[15:12]	);
//SEG7_LUT	u4	(	oSEG4,iDIG[19:16]	);
//SEG7_LUT	u5	(	oSEG5,iDIG[23:20]	);
//SEG7_LUT	u6	(	oSEG6,iDIG[27:24]	);
//SEG7_LUT	u7	(	oSEG7,iDIG[31:28]	);

endmodule