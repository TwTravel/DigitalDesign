// Lookup table used to simplify our pipeline by removing a divide
// Calculates (pixelX - 160)/320 and (pixelY - 120)/240
module pixelRayScaleTable(clk, pixelX, pixelX_minus_160_div_320, pixelY, pixelY_minus_120_div_240);

parameter BusWidth = 0;
parameter DecimalWidth = 0;

input clk;
input [8:0] pixelX, pixelY;
output [BusWidth-1:0] pixelX_minus_160_div_320, pixelY_minus_120_div_240;

reg [15:0] pixelX_minus_160_div_320_16, pixelY_minus_120_div_240_16;

assign pixelX_minus_160_div_320 = {{(BusWidth-DecimalWidth){pixelX_minus_160_div_320_16[15]}}
									,pixelX_minus_160_div_320_16[15:16-DecimalWidth]};
assign pixelY_minus_120_div_240 = {{(BusWidth-DecimalWidth){pixelY_minus_120_div_240_16[15]}}
									,pixelY_minus_120_div_240_16[15:16-DecimalWidth]};

always @(posedge clk)
begin
	case (pixelX)
        9'd0: pixelX_minus_160_div_320_16 <= 16'h8000;
        9'd1: pixelX_minus_160_div_320_16 <= 16'h80cd;
        9'd2: pixelX_minus_160_div_320_16 <= 16'h819a;
        9'd3: pixelX_minus_160_div_320_16 <= 16'h8267;
        9'd4: pixelX_minus_160_div_320_16 <= 16'h8334;
        9'd5: pixelX_minus_160_div_320_16 <= 16'h8400;
        9'd6: pixelX_minus_160_div_320_16 <= 16'h84cd;
        9'd7: pixelX_minus_160_div_320_16 <= 16'h859a;
        9'd8: pixelX_minus_160_div_320_16 <= 16'h8667;
        9'd9: pixelX_minus_160_div_320_16 <= 16'h8734;
        9'd10: pixelX_minus_160_div_320_16 <= 16'h8800;
        9'd11: pixelX_minus_160_div_320_16 <= 16'h88cd;
        9'd12: pixelX_minus_160_div_320_16 <= 16'h899a;
        9'd13: pixelX_minus_160_div_320_16 <= 16'h8a67;
        9'd14: pixelX_minus_160_div_320_16 <= 16'h8b34;
        9'd15: pixelX_minus_160_div_320_16 <= 16'h8c00;
        9'd16: pixelX_minus_160_div_320_16 <= 16'h8ccd;
        9'd17: pixelX_minus_160_div_320_16 <= 16'h8d9a;
        9'd18: pixelX_minus_160_div_320_16 <= 16'h8e67;
        9'd19: pixelX_minus_160_div_320_16 <= 16'h8f34;
        9'd20: pixelX_minus_160_div_320_16 <= 16'h9000;
        9'd21: pixelX_minus_160_div_320_16 <= 16'h90cd;
        9'd22: pixelX_minus_160_div_320_16 <= 16'h919a;
        9'd23: pixelX_minus_160_div_320_16 <= 16'h9267;
        9'd24: pixelX_minus_160_div_320_16 <= 16'h9334;
        9'd25: pixelX_minus_160_div_320_16 <= 16'h9400;
        9'd26: pixelX_minus_160_div_320_16 <= 16'h94cd;
        9'd27: pixelX_minus_160_div_320_16 <= 16'h959a;
        9'd28: pixelX_minus_160_div_320_16 <= 16'h9667;
        9'd29: pixelX_minus_160_div_320_16 <= 16'h9734;
        9'd30: pixelX_minus_160_div_320_16 <= 16'h9800;
        9'd31: pixelX_minus_160_div_320_16 <= 16'h98cd;
        9'd32: pixelX_minus_160_div_320_16 <= 16'h999a;
        9'd33: pixelX_minus_160_div_320_16 <= 16'h9a67;
        9'd34: pixelX_minus_160_div_320_16 <= 16'h9b34;
        9'd35: pixelX_minus_160_div_320_16 <= 16'h9c00;
        9'd36: pixelX_minus_160_div_320_16 <= 16'h9ccd;
        9'd37: pixelX_minus_160_div_320_16 <= 16'h9d9a;
        9'd38: pixelX_minus_160_div_320_16 <= 16'h9e67;
        9'd39: pixelX_minus_160_div_320_16 <= 16'h9f34;
        9'd40: pixelX_minus_160_div_320_16 <= 16'ha000;
        9'd41: pixelX_minus_160_div_320_16 <= 16'ha0cd;
        9'd42: pixelX_minus_160_div_320_16 <= 16'ha19a;
        9'd43: pixelX_minus_160_div_320_16 <= 16'ha267;
        9'd44: pixelX_minus_160_div_320_16 <= 16'ha334;
        9'd45: pixelX_minus_160_div_320_16 <= 16'ha400;
        9'd46: pixelX_minus_160_div_320_16 <= 16'ha4cd;
        9'd47: pixelX_minus_160_div_320_16 <= 16'ha59a;
        9'd48: pixelX_minus_160_div_320_16 <= 16'ha667;
        9'd49: pixelX_minus_160_div_320_16 <= 16'ha734;
        9'd50: pixelX_minus_160_div_320_16 <= 16'ha800;
        9'd51: pixelX_minus_160_div_320_16 <= 16'ha8cd;
        9'd52: pixelX_minus_160_div_320_16 <= 16'ha99a;
        9'd53: pixelX_minus_160_div_320_16 <= 16'haa67;
        9'd54: pixelX_minus_160_div_320_16 <= 16'hab34;
        9'd55: pixelX_minus_160_div_320_16 <= 16'hac00;
        9'd56: pixelX_minus_160_div_320_16 <= 16'haccd;
        9'd57: pixelX_minus_160_div_320_16 <= 16'had9a;
        9'd58: pixelX_minus_160_div_320_16 <= 16'hae67;
        9'd59: pixelX_minus_160_div_320_16 <= 16'haf34;
        9'd60: pixelX_minus_160_div_320_16 <= 16'hb000;
        9'd61: pixelX_minus_160_div_320_16 <= 16'hb0cd;
        9'd62: pixelX_minus_160_div_320_16 <= 16'hb19a;
        9'd63: pixelX_minus_160_div_320_16 <= 16'hb267;
        9'd64: pixelX_minus_160_div_320_16 <= 16'hb334;
        9'd65: pixelX_minus_160_div_320_16 <= 16'hb400;
        9'd66: pixelX_minus_160_div_320_16 <= 16'hb4cd;
        9'd67: pixelX_minus_160_div_320_16 <= 16'hb59a;
        9'd68: pixelX_minus_160_div_320_16 <= 16'hb667;
        9'd69: pixelX_minus_160_div_320_16 <= 16'hb734;
        9'd70: pixelX_minus_160_div_320_16 <= 16'hb800;
        9'd71: pixelX_minus_160_div_320_16 <= 16'hb8cd;
        9'd72: pixelX_minus_160_div_320_16 <= 16'hb99a;
        9'd73: pixelX_minus_160_div_320_16 <= 16'hba67;
        9'd74: pixelX_minus_160_div_320_16 <= 16'hbb34;
        9'd75: pixelX_minus_160_div_320_16 <= 16'hbc00;
        9'd76: pixelX_minus_160_div_320_16 <= 16'hbccd;
        9'd77: pixelX_minus_160_div_320_16 <= 16'hbd9a;
        9'd78: pixelX_minus_160_div_320_16 <= 16'hbe67;
        9'd79: pixelX_minus_160_div_320_16 <= 16'hbf34;
        9'd80: pixelX_minus_160_div_320_16 <= 16'hc000;
        9'd81: pixelX_minus_160_div_320_16 <= 16'hc0cd;
        9'd82: pixelX_minus_160_div_320_16 <= 16'hc19a;
        9'd83: pixelX_minus_160_div_320_16 <= 16'hc267;
        9'd84: pixelX_minus_160_div_320_16 <= 16'hc334;
        9'd85: pixelX_minus_160_div_320_16 <= 16'hc400;
        9'd86: pixelX_minus_160_div_320_16 <= 16'hc4cd;
        9'd87: pixelX_minus_160_div_320_16 <= 16'hc59a;
        9'd88: pixelX_minus_160_div_320_16 <= 16'hc667;
        9'd89: pixelX_minus_160_div_320_16 <= 16'hc734;
        9'd90: pixelX_minus_160_div_320_16 <= 16'hc800;
        9'd91: pixelX_minus_160_div_320_16 <= 16'hc8cd;
        9'd92: pixelX_minus_160_div_320_16 <= 16'hc99a;
        9'd93: pixelX_minus_160_div_320_16 <= 16'hca67;
        9'd94: pixelX_minus_160_div_320_16 <= 16'hcb34;
        9'd95: pixelX_minus_160_div_320_16 <= 16'hcc00;
        9'd96: pixelX_minus_160_div_320_16 <= 16'hcccd;
        9'd97: pixelX_minus_160_div_320_16 <= 16'hcd9a;
        9'd98: pixelX_minus_160_div_320_16 <= 16'hce67;
        9'd99: pixelX_minus_160_div_320_16 <= 16'hcf34;
        9'd100: pixelX_minus_160_div_320_16 <= 16'hd000;
        9'd101: pixelX_minus_160_div_320_16 <= 16'hd0cd;
        9'd102: pixelX_minus_160_div_320_16 <= 16'hd19a;
        9'd103: pixelX_minus_160_div_320_16 <= 16'hd267;
        9'd104: pixelX_minus_160_div_320_16 <= 16'hd334;
        9'd105: pixelX_minus_160_div_320_16 <= 16'hd400;
        9'd106: pixelX_minus_160_div_320_16 <= 16'hd4cd;
        9'd107: pixelX_minus_160_div_320_16 <= 16'hd59a;
        9'd108: pixelX_minus_160_div_320_16 <= 16'hd667;
        9'd109: pixelX_minus_160_div_320_16 <= 16'hd734;
        9'd110: pixelX_minus_160_div_320_16 <= 16'hd800;
        9'd111: pixelX_minus_160_div_320_16 <= 16'hd8cd;
        9'd112: pixelX_minus_160_div_320_16 <= 16'hd99a;
        9'd113: pixelX_minus_160_div_320_16 <= 16'hda67;
        9'd114: pixelX_minus_160_div_320_16 <= 16'hdb34;
        9'd115: pixelX_minus_160_div_320_16 <= 16'hdc00;
        9'd116: pixelX_minus_160_div_320_16 <= 16'hdccd;
        9'd117: pixelX_minus_160_div_320_16 <= 16'hdd9a;
        9'd118: pixelX_minus_160_div_320_16 <= 16'hde67;
        9'd119: pixelX_minus_160_div_320_16 <= 16'hdf34;
        9'd120: pixelX_minus_160_div_320_16 <= 16'he000;
        9'd121: pixelX_minus_160_div_320_16 <= 16'he0cd;
        9'd122: pixelX_minus_160_div_320_16 <= 16'he19a;
        9'd123: pixelX_minus_160_div_320_16 <= 16'he267;
        9'd124: pixelX_minus_160_div_320_16 <= 16'he334;
        9'd125: pixelX_minus_160_div_320_16 <= 16'he400;
        9'd126: pixelX_minus_160_div_320_16 <= 16'he4cd;
        9'd127: pixelX_minus_160_div_320_16 <= 16'he59a;
        9'd128: pixelX_minus_160_div_320_16 <= 16'he667;
        9'd129: pixelX_minus_160_div_320_16 <= 16'he734;
        9'd130: pixelX_minus_160_div_320_16 <= 16'he800;
        9'd131: pixelX_minus_160_div_320_16 <= 16'he8cd;
        9'd132: pixelX_minus_160_div_320_16 <= 16'he99a;
        9'd133: pixelX_minus_160_div_320_16 <= 16'hea67;
        9'd134: pixelX_minus_160_div_320_16 <= 16'heb34;
        9'd135: pixelX_minus_160_div_320_16 <= 16'hec00;
        9'd136: pixelX_minus_160_div_320_16 <= 16'heccd;
        9'd137: pixelX_minus_160_div_320_16 <= 16'hed9a;
        9'd138: pixelX_minus_160_div_320_16 <= 16'hee67;
        9'd139: pixelX_minus_160_div_320_16 <= 16'hef34;
        9'd140: pixelX_minus_160_div_320_16 <= 16'hf000;
        9'd141: pixelX_minus_160_div_320_16 <= 16'hf0cd;
        9'd142: pixelX_minus_160_div_320_16 <= 16'hf19a;
        9'd143: pixelX_minus_160_div_320_16 <= 16'hf267;
        9'd144: pixelX_minus_160_div_320_16 <= 16'hf334;
        9'd145: pixelX_minus_160_div_320_16 <= 16'hf400;
        9'd146: pixelX_minus_160_div_320_16 <= 16'hf4cd;
        9'd147: pixelX_minus_160_div_320_16 <= 16'hf59a;
        9'd148: pixelX_minus_160_div_320_16 <= 16'hf667;
        9'd149: pixelX_minus_160_div_320_16 <= 16'hf734;
        9'd150: pixelX_minus_160_div_320_16 <= 16'hf800;
        9'd151: pixelX_minus_160_div_320_16 <= 16'hf8cd;
        9'd152: pixelX_minus_160_div_320_16 <= 16'hf99a;
        9'd153: pixelX_minus_160_div_320_16 <= 16'hfa67;
        9'd154: pixelX_minus_160_div_320_16 <= 16'hfb34;
        9'd155: pixelX_minus_160_div_320_16 <= 16'hfc00;
        9'd156: pixelX_minus_160_div_320_16 <= 16'hfccd;
        9'd157: pixelX_minus_160_div_320_16 <= 16'hfd9a;
        9'd158: pixelX_minus_160_div_320_16 <= 16'hfe67;
        9'd159: pixelX_minus_160_div_320_16 <= 16'hff34;
        9'd160: pixelX_minus_160_div_320_16 <= 16'h0000;
        9'd161: pixelX_minus_160_div_320_16 <= 16'h00cc;
        9'd162: pixelX_minus_160_div_320_16 <= 16'h0199;
        9'd163: pixelX_minus_160_div_320_16 <= 16'h0266;
        9'd164: pixelX_minus_160_div_320_16 <= 16'h0333;
        9'd165: pixelX_minus_160_div_320_16 <= 16'h0400;
        9'd166: pixelX_minus_160_div_320_16 <= 16'h04cc;
        9'd167: pixelX_minus_160_div_320_16 <= 16'h0599;
        9'd168: pixelX_minus_160_div_320_16 <= 16'h0666;
        9'd169: pixelX_minus_160_div_320_16 <= 16'h0733;
        9'd170: pixelX_minus_160_div_320_16 <= 16'h0800;
        9'd171: pixelX_minus_160_div_320_16 <= 16'h08cc;
        9'd172: pixelX_minus_160_div_320_16 <= 16'h0999;
        9'd173: pixelX_minus_160_div_320_16 <= 16'h0a66;
        9'd174: pixelX_minus_160_div_320_16 <= 16'h0b33;
        9'd175: pixelX_minus_160_div_320_16 <= 16'h0c00;
        9'd176: pixelX_minus_160_div_320_16 <= 16'h0ccc;
        9'd177: pixelX_minus_160_div_320_16 <= 16'h0d99;
        9'd178: pixelX_minus_160_div_320_16 <= 16'h0e66;
        9'd179: pixelX_minus_160_div_320_16 <= 16'h0f33;
        9'd180: pixelX_minus_160_div_320_16 <= 16'h1000;
        9'd181: pixelX_minus_160_div_320_16 <= 16'h10cc;
        9'd182: pixelX_minus_160_div_320_16 <= 16'h1199;
        9'd183: pixelX_minus_160_div_320_16 <= 16'h1266;
        9'd184: pixelX_minus_160_div_320_16 <= 16'h1333;
        9'd185: pixelX_minus_160_div_320_16 <= 16'h1400;
        9'd186: pixelX_minus_160_div_320_16 <= 16'h14cc;
        9'd187: pixelX_minus_160_div_320_16 <= 16'h1599;
        9'd188: pixelX_minus_160_div_320_16 <= 16'h1666;
        9'd189: pixelX_minus_160_div_320_16 <= 16'h1733;
        9'd190: pixelX_minus_160_div_320_16 <= 16'h1800;
        9'd191: pixelX_minus_160_div_320_16 <= 16'h18cc;
        9'd192: pixelX_minus_160_div_320_16 <= 16'h1999;
        9'd193: pixelX_minus_160_div_320_16 <= 16'h1a66;
        9'd194: pixelX_minus_160_div_320_16 <= 16'h1b33;
        9'd195: pixelX_minus_160_div_320_16 <= 16'h1c00;
        9'd196: pixelX_minus_160_div_320_16 <= 16'h1ccc;
        9'd197: pixelX_minus_160_div_320_16 <= 16'h1d99;
        9'd198: pixelX_minus_160_div_320_16 <= 16'h1e66;
        9'd199: pixelX_minus_160_div_320_16 <= 16'h1f33;
        9'd200: pixelX_minus_160_div_320_16 <= 16'h2000;
        9'd201: pixelX_minus_160_div_320_16 <= 16'h20cc;
        9'd202: pixelX_minus_160_div_320_16 <= 16'h2199;
        9'd203: pixelX_minus_160_div_320_16 <= 16'h2266;
        9'd204: pixelX_minus_160_div_320_16 <= 16'h2333;
        9'd205: pixelX_minus_160_div_320_16 <= 16'h2400;
        9'd206: pixelX_minus_160_div_320_16 <= 16'h24cc;
        9'd207: pixelX_minus_160_div_320_16 <= 16'h2599;
        9'd208: pixelX_minus_160_div_320_16 <= 16'h2666;
        9'd209: pixelX_minus_160_div_320_16 <= 16'h2733;
        9'd210: pixelX_minus_160_div_320_16 <= 16'h2800;
        9'd211: pixelX_minus_160_div_320_16 <= 16'h28cc;
        9'd212: pixelX_minus_160_div_320_16 <= 16'h2999;
        9'd213: pixelX_minus_160_div_320_16 <= 16'h2a66;
        9'd214: pixelX_minus_160_div_320_16 <= 16'h2b33;
        9'd215: pixelX_minus_160_div_320_16 <= 16'h2c00;
        9'd216: pixelX_minus_160_div_320_16 <= 16'h2ccc;
        9'd217: pixelX_minus_160_div_320_16 <= 16'h2d99;
        9'd218: pixelX_minus_160_div_320_16 <= 16'h2e66;
        9'd219: pixelX_minus_160_div_320_16 <= 16'h2f33;
        9'd220: pixelX_minus_160_div_320_16 <= 16'h3000;
        9'd221: pixelX_minus_160_div_320_16 <= 16'h30cc;
        9'd222: pixelX_minus_160_div_320_16 <= 16'h3199;
        9'd223: pixelX_minus_160_div_320_16 <= 16'h3266;
        9'd224: pixelX_minus_160_div_320_16 <= 16'h3333;
        9'd225: pixelX_minus_160_div_320_16 <= 16'h3400;
        9'd226: pixelX_minus_160_div_320_16 <= 16'h34cc;
        9'd227: pixelX_minus_160_div_320_16 <= 16'h3599;
        9'd228: pixelX_minus_160_div_320_16 <= 16'h3666;
        9'd229: pixelX_minus_160_div_320_16 <= 16'h3733;
        9'd230: pixelX_minus_160_div_320_16 <= 16'h3800;
        9'd231: pixelX_minus_160_div_320_16 <= 16'h38cc;
        9'd232: pixelX_minus_160_div_320_16 <= 16'h3999;
        9'd233: pixelX_minus_160_div_320_16 <= 16'h3a66;
        9'd234: pixelX_minus_160_div_320_16 <= 16'h3b33;
        9'd235: pixelX_minus_160_div_320_16 <= 16'h3c00;
        9'd236: pixelX_minus_160_div_320_16 <= 16'h3ccc;
        9'd237: pixelX_minus_160_div_320_16 <= 16'h3d99;
        9'd238: pixelX_minus_160_div_320_16 <= 16'h3e66;
        9'd239: pixelX_minus_160_div_320_16 <= 16'h3f33;
        9'd240: pixelX_minus_160_div_320_16 <= 16'h4000;
        9'd241: pixelX_minus_160_div_320_16 <= 16'h40cc;
        9'd242: pixelX_minus_160_div_320_16 <= 16'h4199;
        9'd243: pixelX_minus_160_div_320_16 <= 16'h4266;
        9'd244: pixelX_minus_160_div_320_16 <= 16'h4333;
        9'd245: pixelX_minus_160_div_320_16 <= 16'h4400;
        9'd246: pixelX_minus_160_div_320_16 <= 16'h44cc;
        9'd247: pixelX_minus_160_div_320_16 <= 16'h4599;
        9'd248: pixelX_minus_160_div_320_16 <= 16'h4666;
        9'd249: pixelX_minus_160_div_320_16 <= 16'h4733;
        9'd250: pixelX_minus_160_div_320_16 <= 16'h4800;
        9'd251: pixelX_minus_160_div_320_16 <= 16'h48cc;
        9'd252: pixelX_minus_160_div_320_16 <= 16'h4999;
        9'd253: pixelX_minus_160_div_320_16 <= 16'h4a66;
        9'd254: pixelX_minus_160_div_320_16 <= 16'h4b33;
        9'd255: pixelX_minus_160_div_320_16 <= 16'h4c00;
        9'd256: pixelX_minus_160_div_320_16 <= 16'h4ccc;
        9'd257: pixelX_minus_160_div_320_16 <= 16'h4d99;
        9'd258: pixelX_minus_160_div_320_16 <= 16'h4e66;
        9'd259: pixelX_minus_160_div_320_16 <= 16'h4f33;
        9'd260: pixelX_minus_160_div_320_16 <= 16'h5000;
        9'd261: pixelX_minus_160_div_320_16 <= 16'h50cc;
        9'd262: pixelX_minus_160_div_320_16 <= 16'h5199;
        9'd263: pixelX_minus_160_div_320_16 <= 16'h5266;
        9'd264: pixelX_minus_160_div_320_16 <= 16'h5333;
        9'd265: pixelX_minus_160_div_320_16 <= 16'h5400;
        9'd266: pixelX_minus_160_div_320_16 <= 16'h54cc;
        9'd267: pixelX_minus_160_div_320_16 <= 16'h5599;
        9'd268: pixelX_minus_160_div_320_16 <= 16'h5666;
        9'd269: pixelX_minus_160_div_320_16 <= 16'h5733;
        9'd270: pixelX_minus_160_div_320_16 <= 16'h5800;
        9'd271: pixelX_minus_160_div_320_16 <= 16'h58cc;
        9'd272: pixelX_minus_160_div_320_16 <= 16'h5999;
        9'd273: pixelX_minus_160_div_320_16 <= 16'h5a66;
        9'd274: pixelX_minus_160_div_320_16 <= 16'h5b33;
        9'd275: pixelX_minus_160_div_320_16 <= 16'h5c00;
        9'd276: pixelX_minus_160_div_320_16 <= 16'h5ccc;
        9'd277: pixelX_minus_160_div_320_16 <= 16'h5d99;
        9'd278: pixelX_minus_160_div_320_16 <= 16'h5e66;
        9'd279: pixelX_minus_160_div_320_16 <= 16'h5f33;
        9'd280: pixelX_minus_160_div_320_16 <= 16'h6000;
        9'd281: pixelX_minus_160_div_320_16 <= 16'h60cc;
        9'd282: pixelX_minus_160_div_320_16 <= 16'h6199;
        9'd283: pixelX_minus_160_div_320_16 <= 16'h6266;
        9'd284: pixelX_minus_160_div_320_16 <= 16'h6333;
        9'd285: pixelX_minus_160_div_320_16 <= 16'h6400;
        9'd286: pixelX_minus_160_div_320_16 <= 16'h64cc;
        9'd287: pixelX_minus_160_div_320_16 <= 16'h6599;
        9'd288: pixelX_minus_160_div_320_16 <= 16'h6666;
        9'd289: pixelX_minus_160_div_320_16 <= 16'h6733;
        9'd290: pixelX_minus_160_div_320_16 <= 16'h6800;
        9'd291: pixelX_minus_160_div_320_16 <= 16'h68cc;
        9'd292: pixelX_minus_160_div_320_16 <= 16'h6999;
        9'd293: pixelX_minus_160_div_320_16 <= 16'h6a66;
        9'd294: pixelX_minus_160_div_320_16 <= 16'h6b33;
        9'd295: pixelX_minus_160_div_320_16 <= 16'h6c00;
        9'd296: pixelX_minus_160_div_320_16 <= 16'h6ccc;
        9'd297: pixelX_minus_160_div_320_16 <= 16'h6d99;
        9'd298: pixelX_minus_160_div_320_16 <= 16'h6e66;
        9'd299: pixelX_minus_160_div_320_16 <= 16'h6f33;
        9'd300: pixelX_minus_160_div_320_16 <= 16'h7000;
        9'd301: pixelX_minus_160_div_320_16 <= 16'h70cc;
        9'd302: pixelX_minus_160_div_320_16 <= 16'h7199;
        9'd303: pixelX_minus_160_div_320_16 <= 16'h7266;
        9'd304: pixelX_minus_160_div_320_16 <= 16'h7333;
        9'd305: pixelX_minus_160_div_320_16 <= 16'h7400;
        9'd306: pixelX_minus_160_div_320_16 <= 16'h74cc;
        9'd307: pixelX_minus_160_div_320_16 <= 16'h7599;
        9'd308: pixelX_minus_160_div_320_16 <= 16'h7666;
        9'd309: pixelX_minus_160_div_320_16 <= 16'h7733;
        9'd310: pixelX_minus_160_div_320_16 <= 16'h7800;
        9'd311: pixelX_minus_160_div_320_16 <= 16'h78cc;
        9'd312: pixelX_minus_160_div_320_16 <= 16'h7999;
        9'd313: pixelX_minus_160_div_320_16 <= 16'h7a66;
        9'd314: pixelX_minus_160_div_320_16 <= 16'h7b33;
        9'd315: pixelX_minus_160_div_320_16 <= 16'h7c00;
        9'd316: pixelX_minus_160_div_320_16 <= 16'h7ccc;
        9'd317: pixelX_minus_160_div_320_16 <= 16'h7d99;
        9'd318: pixelX_minus_160_div_320_16 <= 16'h7e66;
        9'd319: pixelX_minus_160_div_320_16 <= 16'h7f33;
		default: pixelX_minus_160_div_320_16 <= 16'h0000;
	endcase

	case (pixelY)
        9'd0: pixelY_minus_120_div_240_16 <= 16'h8000;
        9'd1: pixelY_minus_120_div_240_16 <= 16'h8112;
        9'd2: pixelY_minus_120_div_240_16 <= 16'h8223;
        9'd3: pixelY_minus_120_div_240_16 <= 16'h8334;
        9'd4: pixelY_minus_120_div_240_16 <= 16'h8445;
        9'd5: pixelY_minus_120_div_240_16 <= 16'h8556;
        9'd6: pixelY_minus_120_div_240_16 <= 16'h8667;
        9'd7: pixelY_minus_120_div_240_16 <= 16'h8778;
        9'd8: pixelY_minus_120_div_240_16 <= 16'h8889;
        9'd9: pixelY_minus_120_div_240_16 <= 16'h899a;
        9'd10: pixelY_minus_120_div_240_16 <= 16'h8aab;
        9'd11: pixelY_minus_120_div_240_16 <= 16'h8bbc;
        9'd12: pixelY_minus_120_div_240_16 <= 16'h8ccd;
        9'd13: pixelY_minus_120_div_240_16 <= 16'h8dde;
        9'd14: pixelY_minus_120_div_240_16 <= 16'h8eef;
        9'd15: pixelY_minus_120_div_240_16 <= 16'h9000;
        9'd16: pixelY_minus_120_div_240_16 <= 16'h9112;
        9'd17: pixelY_minus_120_div_240_16 <= 16'h9223;
        9'd18: pixelY_minus_120_div_240_16 <= 16'h9334;
        9'd19: pixelY_minus_120_div_240_16 <= 16'h9445;
        9'd20: pixelY_minus_120_div_240_16 <= 16'h9556;
        9'd21: pixelY_minus_120_div_240_16 <= 16'h9667;
        9'd22: pixelY_minus_120_div_240_16 <= 16'h9778;
        9'd23: pixelY_minus_120_div_240_16 <= 16'h9889;
        9'd24: pixelY_minus_120_div_240_16 <= 16'h999a;
        9'd25: pixelY_minus_120_div_240_16 <= 16'h9aab;
        9'd26: pixelY_minus_120_div_240_16 <= 16'h9bbc;
        9'd27: pixelY_minus_120_div_240_16 <= 16'h9ccd;
        9'd28: pixelY_minus_120_div_240_16 <= 16'h9dde;
        9'd29: pixelY_minus_120_div_240_16 <= 16'h9eef;
        9'd30: pixelY_minus_120_div_240_16 <= 16'ha000;
        9'd31: pixelY_minus_120_div_240_16 <= 16'ha112;
        9'd32: pixelY_minus_120_div_240_16 <= 16'ha223;
        9'd33: pixelY_minus_120_div_240_16 <= 16'ha334;
        9'd34: pixelY_minus_120_div_240_16 <= 16'ha445;
        9'd35: pixelY_minus_120_div_240_16 <= 16'ha556;
        9'd36: pixelY_minus_120_div_240_16 <= 16'ha667;
        9'd37: pixelY_minus_120_div_240_16 <= 16'ha778;
        9'd38: pixelY_minus_120_div_240_16 <= 16'ha889;
        9'd39: pixelY_minus_120_div_240_16 <= 16'ha99a;
        9'd40: pixelY_minus_120_div_240_16 <= 16'haaab;
        9'd41: pixelY_minus_120_div_240_16 <= 16'habbc;
        9'd42: pixelY_minus_120_div_240_16 <= 16'haccd;
        9'd43: pixelY_minus_120_div_240_16 <= 16'hadde;
        9'd44: pixelY_minus_120_div_240_16 <= 16'haeef;
        9'd45: pixelY_minus_120_div_240_16 <= 16'hb000;
        9'd46: pixelY_minus_120_div_240_16 <= 16'hb112;
        9'd47: pixelY_minus_120_div_240_16 <= 16'hb223;
        9'd48: pixelY_minus_120_div_240_16 <= 16'hb334;
        9'd49: pixelY_minus_120_div_240_16 <= 16'hb445;
        9'd50: pixelY_minus_120_div_240_16 <= 16'hb556;
        9'd51: pixelY_minus_120_div_240_16 <= 16'hb667;
        9'd52: pixelY_minus_120_div_240_16 <= 16'hb778;
        9'd53: pixelY_minus_120_div_240_16 <= 16'hb889;
        9'd54: pixelY_minus_120_div_240_16 <= 16'hb99a;
        9'd55: pixelY_minus_120_div_240_16 <= 16'hbaab;
        9'd56: pixelY_minus_120_div_240_16 <= 16'hbbbc;
        9'd57: pixelY_minus_120_div_240_16 <= 16'hbccd;
        9'd58: pixelY_minus_120_div_240_16 <= 16'hbdde;
        9'd59: pixelY_minus_120_div_240_16 <= 16'hbeef;
        9'd60: pixelY_minus_120_div_240_16 <= 16'hc000;
        9'd61: pixelY_minus_120_div_240_16 <= 16'hc112;
        9'd62: pixelY_minus_120_div_240_16 <= 16'hc223;
        9'd63: pixelY_minus_120_div_240_16 <= 16'hc334;
        9'd64: pixelY_minus_120_div_240_16 <= 16'hc445;
        9'd65: pixelY_minus_120_div_240_16 <= 16'hc556;
        9'd66: pixelY_minus_120_div_240_16 <= 16'hc667;
        9'd67: pixelY_minus_120_div_240_16 <= 16'hc778;
        9'd68: pixelY_minus_120_div_240_16 <= 16'hc889;
        9'd69: pixelY_minus_120_div_240_16 <= 16'hc99a;
        9'd70: pixelY_minus_120_div_240_16 <= 16'hcaab;
        9'd71: pixelY_minus_120_div_240_16 <= 16'hcbbc;
        9'd72: pixelY_minus_120_div_240_16 <= 16'hcccd;
        9'd73: pixelY_minus_120_div_240_16 <= 16'hcdde;
        9'd74: pixelY_minus_120_div_240_16 <= 16'hceef;
        9'd75: pixelY_minus_120_div_240_16 <= 16'hd000;
        9'd76: pixelY_minus_120_div_240_16 <= 16'hd112;
        9'd77: pixelY_minus_120_div_240_16 <= 16'hd223;
        9'd78: pixelY_minus_120_div_240_16 <= 16'hd334;
        9'd79: pixelY_minus_120_div_240_16 <= 16'hd445;
        9'd80: pixelY_minus_120_div_240_16 <= 16'hd556;
        9'd81: pixelY_minus_120_div_240_16 <= 16'hd667;
        9'd82: pixelY_minus_120_div_240_16 <= 16'hd778;
        9'd83: pixelY_minus_120_div_240_16 <= 16'hd889;
        9'd84: pixelY_minus_120_div_240_16 <= 16'hd99a;
        9'd85: pixelY_minus_120_div_240_16 <= 16'hdaab;
        9'd86: pixelY_minus_120_div_240_16 <= 16'hdbbc;
        9'd87: pixelY_minus_120_div_240_16 <= 16'hdccd;
        9'd88: pixelY_minus_120_div_240_16 <= 16'hddde;
        9'd89: pixelY_minus_120_div_240_16 <= 16'hdeef;
        9'd90: pixelY_minus_120_div_240_16 <= 16'he000;
        9'd91: pixelY_minus_120_div_240_16 <= 16'he112;
        9'd92: pixelY_minus_120_div_240_16 <= 16'he223;
        9'd93: pixelY_minus_120_div_240_16 <= 16'he334;
        9'd94: pixelY_minus_120_div_240_16 <= 16'he445;
        9'd95: pixelY_minus_120_div_240_16 <= 16'he556;
        9'd96: pixelY_minus_120_div_240_16 <= 16'he667;
        9'd97: pixelY_minus_120_div_240_16 <= 16'he778;
        9'd98: pixelY_minus_120_div_240_16 <= 16'he889;
        9'd99: pixelY_minus_120_div_240_16 <= 16'he99a;
        9'd100: pixelY_minus_120_div_240_16 <= 16'heaab;
        9'd101: pixelY_minus_120_div_240_16 <= 16'hebbc;
        9'd102: pixelY_minus_120_div_240_16 <= 16'heccd;
        9'd103: pixelY_minus_120_div_240_16 <= 16'hedde;
        9'd104: pixelY_minus_120_div_240_16 <= 16'heeef;
        9'd105: pixelY_minus_120_div_240_16 <= 16'hf000;
        9'd106: pixelY_minus_120_div_240_16 <= 16'hf112;
        9'd107: pixelY_minus_120_div_240_16 <= 16'hf223;
        9'd108: pixelY_minus_120_div_240_16 <= 16'hf334;
        9'd109: pixelY_minus_120_div_240_16 <= 16'hf445;
        9'd110: pixelY_minus_120_div_240_16 <= 16'hf556;
        9'd111: pixelY_minus_120_div_240_16 <= 16'hf667;
        9'd112: pixelY_minus_120_div_240_16 <= 16'hf778;
        9'd113: pixelY_minus_120_div_240_16 <= 16'hf889;
        9'd114: pixelY_minus_120_div_240_16 <= 16'hf99a;
        9'd115: pixelY_minus_120_div_240_16 <= 16'hfaab;
        9'd116: pixelY_minus_120_div_240_16 <= 16'hfbbc;
        9'd117: pixelY_minus_120_div_240_16 <= 16'hfccd;
        9'd118: pixelY_minus_120_div_240_16 <= 16'hfdde;
        9'd119: pixelY_minus_120_div_240_16 <= 16'hfeef;
        9'd120: pixelY_minus_120_div_240_16 <= 16'h0000;
        9'd121: pixelY_minus_120_div_240_16 <= 16'h0111;
        9'd122: pixelY_minus_120_div_240_16 <= 16'h0222;
        9'd123: pixelY_minus_120_div_240_16 <= 16'h0333;
        9'd124: pixelY_minus_120_div_240_16 <= 16'h0444;
        9'd125: pixelY_minus_120_div_240_16 <= 16'h0555;
        9'd126: pixelY_minus_120_div_240_16 <= 16'h0666;
        9'd127: pixelY_minus_120_div_240_16 <= 16'h0777;
        9'd128: pixelY_minus_120_div_240_16 <= 16'h0888;
        9'd129: pixelY_minus_120_div_240_16 <= 16'h0999;
        9'd130: pixelY_minus_120_div_240_16 <= 16'h0aaa;
        9'd131: pixelY_minus_120_div_240_16 <= 16'h0bbb;
        9'd132: pixelY_minus_120_div_240_16 <= 16'h0ccc;
        9'd133: pixelY_minus_120_div_240_16 <= 16'h0ddd;
        9'd134: pixelY_minus_120_div_240_16 <= 16'h0eee;
        9'd135: pixelY_minus_120_div_240_16 <= 16'h1000;
        9'd136: pixelY_minus_120_div_240_16 <= 16'h1111;
        9'd137: pixelY_minus_120_div_240_16 <= 16'h1222;
        9'd138: pixelY_minus_120_div_240_16 <= 16'h1333;
        9'd139: pixelY_minus_120_div_240_16 <= 16'h1444;
        9'd140: pixelY_minus_120_div_240_16 <= 16'h1555;
        9'd141: pixelY_minus_120_div_240_16 <= 16'h1666;
        9'd142: pixelY_minus_120_div_240_16 <= 16'h1777;
        9'd143: pixelY_minus_120_div_240_16 <= 16'h1888;
        9'd144: pixelY_minus_120_div_240_16 <= 16'h1999;
        9'd145: pixelY_minus_120_div_240_16 <= 16'h1aaa;
        9'd146: pixelY_minus_120_div_240_16 <= 16'h1bbb;
        9'd147: pixelY_minus_120_div_240_16 <= 16'h1ccc;
        9'd148: pixelY_minus_120_div_240_16 <= 16'h1ddd;
        9'd149: pixelY_minus_120_div_240_16 <= 16'h1eee;
        9'd150: pixelY_minus_120_div_240_16 <= 16'h2000;
        9'd151: pixelY_minus_120_div_240_16 <= 16'h2111;
        9'd152: pixelY_minus_120_div_240_16 <= 16'h2222;
        9'd153: pixelY_minus_120_div_240_16 <= 16'h2333;
        9'd154: pixelY_minus_120_div_240_16 <= 16'h2444;
        9'd155: pixelY_minus_120_div_240_16 <= 16'h2555;
        9'd156: pixelY_minus_120_div_240_16 <= 16'h2666;
        9'd157: pixelY_minus_120_div_240_16 <= 16'h2777;
        9'd158: pixelY_minus_120_div_240_16 <= 16'h2888;
        9'd159: pixelY_minus_120_div_240_16 <= 16'h2999;
        9'd160: pixelY_minus_120_div_240_16 <= 16'h2aaa;
        9'd161: pixelY_minus_120_div_240_16 <= 16'h2bbb;
        9'd162: pixelY_minus_120_div_240_16 <= 16'h2ccc;
        9'd163: pixelY_minus_120_div_240_16 <= 16'h2ddd;
        9'd164: pixelY_minus_120_div_240_16 <= 16'h2eee;
        9'd165: pixelY_minus_120_div_240_16 <= 16'h3000;
        9'd166: pixelY_minus_120_div_240_16 <= 16'h3111;
        9'd167: pixelY_minus_120_div_240_16 <= 16'h3222;
        9'd168: pixelY_minus_120_div_240_16 <= 16'h3333;
        9'd169: pixelY_minus_120_div_240_16 <= 16'h3444;
        9'd170: pixelY_minus_120_div_240_16 <= 16'h3555;
        9'd171: pixelY_minus_120_div_240_16 <= 16'h3666;
        9'd172: pixelY_minus_120_div_240_16 <= 16'h3777;
        9'd173: pixelY_minus_120_div_240_16 <= 16'h3888;
        9'd174: pixelY_minus_120_div_240_16 <= 16'h3999;
        9'd175: pixelY_minus_120_div_240_16 <= 16'h3aaa;
        9'd176: pixelY_minus_120_div_240_16 <= 16'h3bbb;
        9'd177: pixelY_minus_120_div_240_16 <= 16'h3ccc;
        9'd178: pixelY_minus_120_div_240_16 <= 16'h3ddd;
        9'd179: pixelY_minus_120_div_240_16 <= 16'h3eee;
        9'd180: pixelY_minus_120_div_240_16 <= 16'h4000;
        9'd181: pixelY_minus_120_div_240_16 <= 16'h4111;
        9'd182: pixelY_minus_120_div_240_16 <= 16'h4222;
        9'd183: pixelY_minus_120_div_240_16 <= 16'h4333;
        9'd184: pixelY_minus_120_div_240_16 <= 16'h4444;
        9'd185: pixelY_minus_120_div_240_16 <= 16'h4555;
        9'd186: pixelY_minus_120_div_240_16 <= 16'h4666;
        9'd187: pixelY_minus_120_div_240_16 <= 16'h4777;
        9'd188: pixelY_minus_120_div_240_16 <= 16'h4888;
        9'd189: pixelY_minus_120_div_240_16 <= 16'h4999;
        9'd190: pixelY_minus_120_div_240_16 <= 16'h4aaa;
        9'd191: pixelY_minus_120_div_240_16 <= 16'h4bbb;
        9'd192: pixelY_minus_120_div_240_16 <= 16'h4ccc;
        9'd193: pixelY_minus_120_div_240_16 <= 16'h4ddd;
        9'd194: pixelY_minus_120_div_240_16 <= 16'h4eee;
        9'd195: pixelY_minus_120_div_240_16 <= 16'h5000;
        9'd196: pixelY_minus_120_div_240_16 <= 16'h5111;
        9'd197: pixelY_minus_120_div_240_16 <= 16'h5222;
        9'd198: pixelY_minus_120_div_240_16 <= 16'h5333;
        9'd199: pixelY_minus_120_div_240_16 <= 16'h5444;
        9'd200: pixelY_minus_120_div_240_16 <= 16'h5555;
        9'd201: pixelY_minus_120_div_240_16 <= 16'h5666;
        9'd202: pixelY_minus_120_div_240_16 <= 16'h5777;
        9'd203: pixelY_minus_120_div_240_16 <= 16'h5888;
        9'd204: pixelY_minus_120_div_240_16 <= 16'h5999;
        9'd205: pixelY_minus_120_div_240_16 <= 16'h5aaa;
        9'd206: pixelY_minus_120_div_240_16 <= 16'h5bbb;
        9'd207: pixelY_minus_120_div_240_16 <= 16'h5ccc;
        9'd208: pixelY_minus_120_div_240_16 <= 16'h5ddd;
        9'd209: pixelY_minus_120_div_240_16 <= 16'h5eee;
        9'd210: pixelY_minus_120_div_240_16 <= 16'h6000;
        9'd211: pixelY_minus_120_div_240_16 <= 16'h6111;
        9'd212: pixelY_minus_120_div_240_16 <= 16'h6222;
        9'd213: pixelY_minus_120_div_240_16 <= 16'h6333;
        9'd214: pixelY_minus_120_div_240_16 <= 16'h6444;
        9'd215: pixelY_minus_120_div_240_16 <= 16'h6555;
        9'd216: pixelY_minus_120_div_240_16 <= 16'h6666;
        9'd217: pixelY_minus_120_div_240_16 <= 16'h6777;
        9'd218: pixelY_minus_120_div_240_16 <= 16'h6888;
        9'd219: pixelY_minus_120_div_240_16 <= 16'h6999;
        9'd220: pixelY_minus_120_div_240_16 <= 16'h6aaa;
        9'd221: pixelY_minus_120_div_240_16 <= 16'h6bbb;
        9'd222: pixelY_minus_120_div_240_16 <= 16'h6ccc;
        9'd223: pixelY_minus_120_div_240_16 <= 16'h6ddd;
        9'd224: pixelY_minus_120_div_240_16 <= 16'h6eee;
        9'd225: pixelY_minus_120_div_240_16 <= 16'h7000;
        9'd226: pixelY_minus_120_div_240_16 <= 16'h7111;
        9'd227: pixelY_minus_120_div_240_16 <= 16'h7222;
        9'd228: pixelY_minus_120_div_240_16 <= 16'h7333;
        9'd229: pixelY_minus_120_div_240_16 <= 16'h7444;
        9'd230: pixelY_minus_120_div_240_16 <= 16'h7555;
        9'd231: pixelY_minus_120_div_240_16 <= 16'h7666;
        9'd232: pixelY_minus_120_div_240_16 <= 16'h7777;
        9'd233: pixelY_minus_120_div_240_16 <= 16'h7888;
        9'd234: pixelY_minus_120_div_240_16 <= 16'h7999;
        9'd235: pixelY_minus_120_div_240_16 <= 16'h7aaa;
        9'd236: pixelY_minus_120_div_240_16 <= 16'h7bbb;
        9'd237: pixelY_minus_120_div_240_16 <= 16'h7ccc;
        9'd238: pixelY_minus_120_div_240_16 <= 16'h7ddd;
        9'd239: pixelY_minus_120_div_240_16 <= 16'h7eee;
		default: pixelY_minus_120_div_240_16 <= 16'h0000;
	endcase				

end


endmodule