/****************************************************************
 * Skyler Schneider ss868                                       *
 * ECE 5760 Final Project                                       *
 * Sand Game                                                    *
 ****************************************************************/

// Produces yes/no answer whether a pixel offset (Xdist, Ydist)
// from the center of a circle is actually within that circle.
module CircleROM (
    input             iCLK,  // Clock signal for reading
    input      [11:0] iAddr, // {CircleSize, Xdist, Ydist}
    output reg        oData  // Pixel value - yes/no answer
);
    
    always @(posedge iCLK) begin
        case(iAddr)
            12'h000: oData <= 1'b1;
            12'h001: oData <= 1'b0;
            12'h002: oData <= 1'b0;
            12'h003: oData <= 1'b0;
            12'h004: oData <= 1'b0;
            12'h005: oData <= 1'b0;
            12'h006: oData <= 1'b0;
            12'h007: oData <= 1'b0;
            12'h008: oData <= 1'b0;
            12'h009: oData <= 1'b0;
            12'h00a: oData <= 1'b0;
            12'h00b: oData <= 1'b0;
            12'h00c: oData <= 1'b0;
            12'h00d: oData <= 1'b0;
            12'h00e: oData <= 1'b0;
            12'h00f: oData <= 1'b0;
            12'h010: oData <= 1'b0;
            12'h011: oData <= 1'b0;
            12'h012: oData <= 1'b0;
            12'h013: oData <= 1'b0;
            12'h014: oData <= 1'b0;
            12'h015: oData <= 1'b0;
            12'h016: oData <= 1'b0;
            12'h017: oData <= 1'b0;
            12'h018: oData <= 1'b0;
            12'h019: oData <= 1'b0;
            12'h01a: oData <= 1'b0;
            12'h01b: oData <= 1'b0;
            12'h01c: oData <= 1'b0;
            12'h01d: oData <= 1'b0;
            12'h01e: oData <= 1'b0;
            12'h01f: oData <= 1'b0;
            12'h020: oData <= 1'b0;
            12'h021: oData <= 1'b0;
            12'h022: oData <= 1'b0;
            12'h023: oData <= 1'b0;
            12'h024: oData <= 1'b0;
            12'h025: oData <= 1'b0;
            12'h026: oData <= 1'b0;
            12'h027: oData <= 1'b0;
            12'h028: oData <= 1'b0;
            12'h029: oData <= 1'b0;
            12'h02a: oData <= 1'b0;
            12'h02b: oData <= 1'b0;
            12'h02c: oData <= 1'b0;
            12'h02d: oData <= 1'b0;
            12'h02e: oData <= 1'b0;
            12'h02f: oData <= 1'b0;
            12'h030: oData <= 1'b0;
            12'h031: oData <= 1'b0;
            12'h032: oData <= 1'b0;
            12'h033: oData <= 1'b0;
            12'h034: oData <= 1'b0;
            12'h035: oData <= 1'b0;
            12'h036: oData <= 1'b0;
            12'h037: oData <= 1'b0;
            12'h038: oData <= 1'b0;
            12'h039: oData <= 1'b0;
            12'h03a: oData <= 1'b0;
            12'h03b: oData <= 1'b0;
            12'h03c: oData <= 1'b0;
            12'h03d: oData <= 1'b0;
            12'h03e: oData <= 1'b0;
            12'h03f: oData <= 1'b0;
            12'h040: oData <= 1'b0;
            12'h041: oData <= 1'b0;
            12'h042: oData <= 1'b0;
            12'h043: oData <= 1'b0;
            12'h044: oData <= 1'b0;
            12'h045: oData <= 1'b0;
            12'h046: oData <= 1'b0;
            12'h047: oData <= 1'b0;
            12'h048: oData <= 1'b0;
            12'h049: oData <= 1'b0;
            12'h04a: oData <= 1'b0;
            12'h04b: oData <= 1'b0;
            12'h04c: oData <= 1'b0;
            12'h04d: oData <= 1'b0;
            12'h04e: oData <= 1'b0;
            12'h04f: oData <= 1'b0;
            12'h050: oData <= 1'b0;
            12'h051: oData <= 1'b0;
            12'h052: oData <= 1'b0;
            12'h053: oData <= 1'b0;
            12'h054: oData <= 1'b0;
            12'h055: oData <= 1'b0;
            12'h056: oData <= 1'b0;
            12'h057: oData <= 1'b0;
            12'h058: oData <= 1'b0;
            12'h059: oData <= 1'b0;
            12'h05a: oData <= 1'b0;
            12'h05b: oData <= 1'b0;
            12'h05c: oData <= 1'b0;
            12'h05d: oData <= 1'b0;
            12'h05e: oData <= 1'b0;
            12'h05f: oData <= 1'b0;
            12'h060: oData <= 1'b0;
            12'h061: oData <= 1'b0;
            12'h062: oData <= 1'b0;
            12'h063: oData <= 1'b0;
            12'h064: oData <= 1'b0;
            12'h065: oData <= 1'b0;
            12'h066: oData <= 1'b0;
            12'h067: oData <= 1'b0;
            12'h068: oData <= 1'b0;
            12'h069: oData <= 1'b0;
            12'h06a: oData <= 1'b0;
            12'h06b: oData <= 1'b0;
            12'h06c: oData <= 1'b0;
            12'h06d: oData <= 1'b0;
            12'h06e: oData <= 1'b0;
            12'h06f: oData <= 1'b0;
            12'h070: oData <= 1'b0;
            12'h071: oData <= 1'b0;
            12'h072: oData <= 1'b0;
            12'h073: oData <= 1'b0;
            12'h074: oData <= 1'b0;
            12'h075: oData <= 1'b0;
            12'h076: oData <= 1'b0;
            12'h077: oData <= 1'b0;
            12'h078: oData <= 1'b0;
            12'h079: oData <= 1'b0;
            12'h07a: oData <= 1'b0;
            12'h07b: oData <= 1'b0;
            12'h07c: oData <= 1'b0;
            12'h07d: oData <= 1'b0;
            12'h07e: oData <= 1'b0;
            12'h07f: oData <= 1'b0;
            12'h080: oData <= 1'b0;
            12'h081: oData <= 1'b0;
            12'h082: oData <= 1'b0;
            12'h083: oData <= 1'b0;
            12'h084: oData <= 1'b0;
            12'h085: oData <= 1'b0;
            12'h086: oData <= 1'b0;
            12'h087: oData <= 1'b0;
            12'h088: oData <= 1'b0;
            12'h089: oData <= 1'b0;
            12'h08a: oData <= 1'b0;
            12'h08b: oData <= 1'b0;
            12'h08c: oData <= 1'b0;
            12'h08d: oData <= 1'b0;
            12'h08e: oData <= 1'b0;
            12'h08f: oData <= 1'b0;
            12'h090: oData <= 1'b0;
            12'h091: oData <= 1'b0;
            12'h092: oData <= 1'b0;
            12'h093: oData <= 1'b0;
            12'h094: oData <= 1'b0;
            12'h095: oData <= 1'b0;
            12'h096: oData <= 1'b0;
            12'h097: oData <= 1'b0;
            12'h098: oData <= 1'b0;
            12'h099: oData <= 1'b0;
            12'h09a: oData <= 1'b0;
            12'h09b: oData <= 1'b0;
            12'h09c: oData <= 1'b0;
            12'h09d: oData <= 1'b0;
            12'h09e: oData <= 1'b0;
            12'h09f: oData <= 1'b0;
            12'h0a0: oData <= 1'b0;
            12'h0a1: oData <= 1'b0;
            12'h0a2: oData <= 1'b0;
            12'h0a3: oData <= 1'b0;
            12'h0a4: oData <= 1'b0;
            12'h0a5: oData <= 1'b0;
            12'h0a6: oData <= 1'b0;
            12'h0a7: oData <= 1'b0;
            12'h0a8: oData <= 1'b0;
            12'h0a9: oData <= 1'b0;
            12'h0aa: oData <= 1'b0;
            12'h0ab: oData <= 1'b0;
            12'h0ac: oData <= 1'b0;
            12'h0ad: oData <= 1'b0;
            12'h0ae: oData <= 1'b0;
            12'h0af: oData <= 1'b0;
            12'h0b0: oData <= 1'b0;
            12'h0b1: oData <= 1'b0;
            12'h0b2: oData <= 1'b0;
            12'h0b3: oData <= 1'b0;
            12'h0b4: oData <= 1'b0;
            12'h0b5: oData <= 1'b0;
            12'h0b6: oData <= 1'b0;
            12'h0b7: oData <= 1'b0;
            12'h0b8: oData <= 1'b0;
            12'h0b9: oData <= 1'b0;
            12'h0ba: oData <= 1'b0;
            12'h0bb: oData <= 1'b0;
            12'h0bc: oData <= 1'b0;
            12'h0bd: oData <= 1'b0;
            12'h0be: oData <= 1'b0;
            12'h0bf: oData <= 1'b0;
            12'h0c0: oData <= 1'b0;
            12'h0c1: oData <= 1'b0;
            12'h0c2: oData <= 1'b0;
            12'h0c3: oData <= 1'b0;
            12'h0c4: oData <= 1'b0;
            12'h0c5: oData <= 1'b0;
            12'h0c6: oData <= 1'b0;
            12'h0c7: oData <= 1'b0;
            12'h0c8: oData <= 1'b0;
            12'h0c9: oData <= 1'b0;
            12'h0ca: oData <= 1'b0;
            12'h0cb: oData <= 1'b0;
            12'h0cc: oData <= 1'b0;
            12'h0cd: oData <= 1'b0;
            12'h0ce: oData <= 1'b0;
            12'h0cf: oData <= 1'b0;
            12'h0d0: oData <= 1'b0;
            12'h0d1: oData <= 1'b0;
            12'h0d2: oData <= 1'b0;
            12'h0d3: oData <= 1'b0;
            12'h0d4: oData <= 1'b0;
            12'h0d5: oData <= 1'b0;
            12'h0d6: oData <= 1'b0;
            12'h0d7: oData <= 1'b0;
            12'h0d8: oData <= 1'b0;
            12'h0d9: oData <= 1'b0;
            12'h0da: oData <= 1'b0;
            12'h0db: oData <= 1'b0;
            12'h0dc: oData <= 1'b0;
            12'h0dd: oData <= 1'b0;
            12'h0de: oData <= 1'b0;
            12'h0df: oData <= 1'b0;
            12'h0e0: oData <= 1'b0;
            12'h0e1: oData <= 1'b0;
            12'h0e2: oData <= 1'b0;
            12'h0e3: oData <= 1'b0;
            12'h0e4: oData <= 1'b0;
            12'h0e5: oData <= 1'b0;
            12'h0e6: oData <= 1'b0;
            12'h0e7: oData <= 1'b0;
            12'h0e8: oData <= 1'b0;
            12'h0e9: oData <= 1'b0;
            12'h0ea: oData <= 1'b0;
            12'h0eb: oData <= 1'b0;
            12'h0ec: oData <= 1'b0;
            12'h0ed: oData <= 1'b0;
            12'h0ee: oData <= 1'b0;
            12'h0ef: oData <= 1'b0;
            12'h0f0: oData <= 1'b0;
            12'h0f1: oData <= 1'b0;
            12'h0f2: oData <= 1'b0;
            12'h0f3: oData <= 1'b0;
            12'h0f4: oData <= 1'b0;
            12'h0f5: oData <= 1'b0;
            12'h0f6: oData <= 1'b0;
            12'h0f7: oData <= 1'b0;
            12'h0f8: oData <= 1'b0;
            12'h0f9: oData <= 1'b0;
            12'h0fa: oData <= 1'b0;
            12'h0fb: oData <= 1'b0;
            12'h0fc: oData <= 1'b0;
            12'h0fd: oData <= 1'b0;
            12'h0fe: oData <= 1'b0;
            12'h0ff: oData <= 1'b0;
            12'h100: oData <= 1'b1;
            12'h101: oData <= 1'b1;
            12'h102: oData <= 1'b0;
            12'h103: oData <= 1'b0;
            12'h104: oData <= 1'b0;
            12'h105: oData <= 1'b0;
            12'h106: oData <= 1'b0;
            12'h107: oData <= 1'b0;
            12'h108: oData <= 1'b0;
            12'h109: oData <= 1'b0;
            12'h10a: oData <= 1'b0;
            12'h10b: oData <= 1'b0;
            12'h10c: oData <= 1'b0;
            12'h10d: oData <= 1'b0;
            12'h10e: oData <= 1'b0;
            12'h10f: oData <= 1'b0;
            12'h110: oData <= 1'b1;
            12'h111: oData <= 1'b0;
            12'h112: oData <= 1'b0;
            12'h113: oData <= 1'b0;
            12'h114: oData <= 1'b0;
            12'h115: oData <= 1'b0;
            12'h116: oData <= 1'b0;
            12'h117: oData <= 1'b0;
            12'h118: oData <= 1'b0;
            12'h119: oData <= 1'b0;
            12'h11a: oData <= 1'b0;
            12'h11b: oData <= 1'b0;
            12'h11c: oData <= 1'b0;
            12'h11d: oData <= 1'b0;
            12'h11e: oData <= 1'b0;
            12'h11f: oData <= 1'b0;
            12'h120: oData <= 1'b0;
            12'h121: oData <= 1'b0;
            12'h122: oData <= 1'b0;
            12'h123: oData <= 1'b0;
            12'h124: oData <= 1'b0;
            12'h125: oData <= 1'b0;
            12'h126: oData <= 1'b0;
            12'h127: oData <= 1'b0;
            12'h128: oData <= 1'b0;
            12'h129: oData <= 1'b0;
            12'h12a: oData <= 1'b0;
            12'h12b: oData <= 1'b0;
            12'h12c: oData <= 1'b0;
            12'h12d: oData <= 1'b0;
            12'h12e: oData <= 1'b0;
            12'h12f: oData <= 1'b0;
            12'h130: oData <= 1'b0;
            12'h131: oData <= 1'b0;
            12'h132: oData <= 1'b0;
            12'h133: oData <= 1'b0;
            12'h134: oData <= 1'b0;
            12'h135: oData <= 1'b0;
            12'h136: oData <= 1'b0;
            12'h137: oData <= 1'b0;
            12'h138: oData <= 1'b0;
            12'h139: oData <= 1'b0;
            12'h13a: oData <= 1'b0;
            12'h13b: oData <= 1'b0;
            12'h13c: oData <= 1'b0;
            12'h13d: oData <= 1'b0;
            12'h13e: oData <= 1'b0;
            12'h13f: oData <= 1'b0;
            12'h140: oData <= 1'b0;
            12'h141: oData <= 1'b0;
            12'h142: oData <= 1'b0;
            12'h143: oData <= 1'b0;
            12'h144: oData <= 1'b0;
            12'h145: oData <= 1'b0;
            12'h146: oData <= 1'b0;
            12'h147: oData <= 1'b0;
            12'h148: oData <= 1'b0;
            12'h149: oData <= 1'b0;
            12'h14a: oData <= 1'b0;
            12'h14b: oData <= 1'b0;
            12'h14c: oData <= 1'b0;
            12'h14d: oData <= 1'b0;
            12'h14e: oData <= 1'b0;
            12'h14f: oData <= 1'b0;
            12'h150: oData <= 1'b0;
            12'h151: oData <= 1'b0;
            12'h152: oData <= 1'b0;
            12'h153: oData <= 1'b0;
            12'h154: oData <= 1'b0;
            12'h155: oData <= 1'b0;
            12'h156: oData <= 1'b0;
            12'h157: oData <= 1'b0;
            12'h158: oData <= 1'b0;
            12'h159: oData <= 1'b0;
            12'h15a: oData <= 1'b0;
            12'h15b: oData <= 1'b0;
            12'h15c: oData <= 1'b0;
            12'h15d: oData <= 1'b0;
            12'h15e: oData <= 1'b0;
            12'h15f: oData <= 1'b0;
            12'h160: oData <= 1'b0;
            12'h161: oData <= 1'b0;
            12'h162: oData <= 1'b0;
            12'h163: oData <= 1'b0;
            12'h164: oData <= 1'b0;
            12'h165: oData <= 1'b0;
            12'h166: oData <= 1'b0;
            12'h167: oData <= 1'b0;
            12'h168: oData <= 1'b0;
            12'h169: oData <= 1'b0;
            12'h16a: oData <= 1'b0;
            12'h16b: oData <= 1'b0;
            12'h16c: oData <= 1'b0;
            12'h16d: oData <= 1'b0;
            12'h16e: oData <= 1'b0;
            12'h16f: oData <= 1'b0;
            12'h170: oData <= 1'b0;
            12'h171: oData <= 1'b0;
            12'h172: oData <= 1'b0;
            12'h173: oData <= 1'b0;
            12'h174: oData <= 1'b0;
            12'h175: oData <= 1'b0;
            12'h176: oData <= 1'b0;
            12'h177: oData <= 1'b0;
            12'h178: oData <= 1'b0;
            12'h179: oData <= 1'b0;
            12'h17a: oData <= 1'b0;
            12'h17b: oData <= 1'b0;
            12'h17c: oData <= 1'b0;
            12'h17d: oData <= 1'b0;
            12'h17e: oData <= 1'b0;
            12'h17f: oData <= 1'b0;
            12'h180: oData <= 1'b0;
            12'h181: oData <= 1'b0;
            12'h182: oData <= 1'b0;
            12'h183: oData <= 1'b0;
            12'h184: oData <= 1'b0;
            12'h185: oData <= 1'b0;
            12'h186: oData <= 1'b0;
            12'h187: oData <= 1'b0;
            12'h188: oData <= 1'b0;
            12'h189: oData <= 1'b0;
            12'h18a: oData <= 1'b0;
            12'h18b: oData <= 1'b0;
            12'h18c: oData <= 1'b0;
            12'h18d: oData <= 1'b0;
            12'h18e: oData <= 1'b0;
            12'h18f: oData <= 1'b0;
            12'h190: oData <= 1'b0;
            12'h191: oData <= 1'b0;
            12'h192: oData <= 1'b0;
            12'h193: oData <= 1'b0;
            12'h194: oData <= 1'b0;
            12'h195: oData <= 1'b0;
            12'h196: oData <= 1'b0;
            12'h197: oData <= 1'b0;
            12'h198: oData <= 1'b0;
            12'h199: oData <= 1'b0;
            12'h19a: oData <= 1'b0;
            12'h19b: oData <= 1'b0;
            12'h19c: oData <= 1'b0;
            12'h19d: oData <= 1'b0;
            12'h19e: oData <= 1'b0;
            12'h19f: oData <= 1'b0;
            12'h1a0: oData <= 1'b0;
            12'h1a1: oData <= 1'b0;
            12'h1a2: oData <= 1'b0;
            12'h1a3: oData <= 1'b0;
            12'h1a4: oData <= 1'b0;
            12'h1a5: oData <= 1'b0;
            12'h1a6: oData <= 1'b0;
            12'h1a7: oData <= 1'b0;
            12'h1a8: oData <= 1'b0;
            12'h1a9: oData <= 1'b0;
            12'h1aa: oData <= 1'b0;
            12'h1ab: oData <= 1'b0;
            12'h1ac: oData <= 1'b0;
            12'h1ad: oData <= 1'b0;
            12'h1ae: oData <= 1'b0;
            12'h1af: oData <= 1'b0;
            12'h1b0: oData <= 1'b0;
            12'h1b1: oData <= 1'b0;
            12'h1b2: oData <= 1'b0;
            12'h1b3: oData <= 1'b0;
            12'h1b4: oData <= 1'b0;
            12'h1b5: oData <= 1'b0;
            12'h1b6: oData <= 1'b0;
            12'h1b7: oData <= 1'b0;
            12'h1b8: oData <= 1'b0;
            12'h1b9: oData <= 1'b0;
            12'h1ba: oData <= 1'b0;
            12'h1bb: oData <= 1'b0;
            12'h1bc: oData <= 1'b0;
            12'h1bd: oData <= 1'b0;
            12'h1be: oData <= 1'b0;
            12'h1bf: oData <= 1'b0;
            12'h1c0: oData <= 1'b0;
            12'h1c1: oData <= 1'b0;
            12'h1c2: oData <= 1'b0;
            12'h1c3: oData <= 1'b0;
            12'h1c4: oData <= 1'b0;
            12'h1c5: oData <= 1'b0;
            12'h1c6: oData <= 1'b0;
            12'h1c7: oData <= 1'b0;
            12'h1c8: oData <= 1'b0;
            12'h1c9: oData <= 1'b0;
            12'h1ca: oData <= 1'b0;
            12'h1cb: oData <= 1'b0;
            12'h1cc: oData <= 1'b0;
            12'h1cd: oData <= 1'b0;
            12'h1ce: oData <= 1'b0;
            12'h1cf: oData <= 1'b0;
            12'h1d0: oData <= 1'b0;
            12'h1d1: oData <= 1'b0;
            12'h1d2: oData <= 1'b0;
            12'h1d3: oData <= 1'b0;
            12'h1d4: oData <= 1'b0;
            12'h1d5: oData <= 1'b0;
            12'h1d6: oData <= 1'b0;
            12'h1d7: oData <= 1'b0;
            12'h1d8: oData <= 1'b0;
            12'h1d9: oData <= 1'b0;
            12'h1da: oData <= 1'b0;
            12'h1db: oData <= 1'b0;
            12'h1dc: oData <= 1'b0;
            12'h1dd: oData <= 1'b0;
            12'h1de: oData <= 1'b0;
            12'h1df: oData <= 1'b0;
            12'h1e0: oData <= 1'b0;
            12'h1e1: oData <= 1'b0;
            12'h1e2: oData <= 1'b0;
            12'h1e3: oData <= 1'b0;
            12'h1e4: oData <= 1'b0;
            12'h1e5: oData <= 1'b0;
            12'h1e6: oData <= 1'b0;
            12'h1e7: oData <= 1'b0;
            12'h1e8: oData <= 1'b0;
            12'h1e9: oData <= 1'b0;
            12'h1ea: oData <= 1'b0;
            12'h1eb: oData <= 1'b0;
            12'h1ec: oData <= 1'b0;
            12'h1ed: oData <= 1'b0;
            12'h1ee: oData <= 1'b0;
            12'h1ef: oData <= 1'b0;
            12'h1f0: oData <= 1'b0;
            12'h1f1: oData <= 1'b0;
            12'h1f2: oData <= 1'b0;
            12'h1f3: oData <= 1'b0;
            12'h1f4: oData <= 1'b0;
            12'h1f5: oData <= 1'b0;
            12'h1f6: oData <= 1'b0;
            12'h1f7: oData <= 1'b0;
            12'h1f8: oData <= 1'b0;
            12'h1f9: oData <= 1'b0;
            12'h1fa: oData <= 1'b0;
            12'h1fb: oData <= 1'b0;
            12'h1fc: oData <= 1'b0;
            12'h1fd: oData <= 1'b0;
            12'h1fe: oData <= 1'b0;
            12'h1ff: oData <= 1'b0;
            12'h200: oData <= 1'b1;
            12'h201: oData <= 1'b1;
            12'h202: oData <= 1'b1;
            12'h203: oData <= 1'b0;
            12'h204: oData <= 1'b0;
            12'h205: oData <= 1'b0;
            12'h206: oData <= 1'b0;
            12'h207: oData <= 1'b0;
            12'h208: oData <= 1'b0;
            12'h209: oData <= 1'b0;
            12'h20a: oData <= 1'b0;
            12'h20b: oData <= 1'b0;
            12'h20c: oData <= 1'b0;
            12'h20d: oData <= 1'b0;
            12'h20e: oData <= 1'b0;
            12'h20f: oData <= 1'b0;
            12'h210: oData <= 1'b1;
            12'h211: oData <= 1'b1;
            12'h212: oData <= 1'b1;
            12'h213: oData <= 1'b0;
            12'h214: oData <= 1'b0;
            12'h215: oData <= 1'b0;
            12'h216: oData <= 1'b0;
            12'h217: oData <= 1'b0;
            12'h218: oData <= 1'b0;
            12'h219: oData <= 1'b0;
            12'h21a: oData <= 1'b0;
            12'h21b: oData <= 1'b0;
            12'h21c: oData <= 1'b0;
            12'h21d: oData <= 1'b0;
            12'h21e: oData <= 1'b0;
            12'h21f: oData <= 1'b0;
            12'h220: oData <= 1'b1;
            12'h221: oData <= 1'b1;
            12'h222: oData <= 1'b0;
            12'h223: oData <= 1'b0;
            12'h224: oData <= 1'b0;
            12'h225: oData <= 1'b0;
            12'h226: oData <= 1'b0;
            12'h227: oData <= 1'b0;
            12'h228: oData <= 1'b0;
            12'h229: oData <= 1'b0;
            12'h22a: oData <= 1'b0;
            12'h22b: oData <= 1'b0;
            12'h22c: oData <= 1'b0;
            12'h22d: oData <= 1'b0;
            12'h22e: oData <= 1'b0;
            12'h22f: oData <= 1'b0;
            12'h230: oData <= 1'b0;
            12'h231: oData <= 1'b0;
            12'h232: oData <= 1'b0;
            12'h233: oData <= 1'b0;
            12'h234: oData <= 1'b0;
            12'h235: oData <= 1'b0;
            12'h236: oData <= 1'b0;
            12'h237: oData <= 1'b0;
            12'h238: oData <= 1'b0;
            12'h239: oData <= 1'b0;
            12'h23a: oData <= 1'b0;
            12'h23b: oData <= 1'b0;
            12'h23c: oData <= 1'b0;
            12'h23d: oData <= 1'b0;
            12'h23e: oData <= 1'b0;
            12'h23f: oData <= 1'b0;
            12'h240: oData <= 1'b0;
            12'h241: oData <= 1'b0;
            12'h242: oData <= 1'b0;
            12'h243: oData <= 1'b0;
            12'h244: oData <= 1'b0;
            12'h245: oData <= 1'b0;
            12'h246: oData <= 1'b0;
            12'h247: oData <= 1'b0;
            12'h248: oData <= 1'b0;
            12'h249: oData <= 1'b0;
            12'h24a: oData <= 1'b0;
            12'h24b: oData <= 1'b0;
            12'h24c: oData <= 1'b0;
            12'h24d: oData <= 1'b0;
            12'h24e: oData <= 1'b0;
            12'h24f: oData <= 1'b0;
            12'h250: oData <= 1'b0;
            12'h251: oData <= 1'b0;
            12'h252: oData <= 1'b0;
            12'h253: oData <= 1'b0;
            12'h254: oData <= 1'b0;
            12'h255: oData <= 1'b0;
            12'h256: oData <= 1'b0;
            12'h257: oData <= 1'b0;
            12'h258: oData <= 1'b0;
            12'h259: oData <= 1'b0;
            12'h25a: oData <= 1'b0;
            12'h25b: oData <= 1'b0;
            12'h25c: oData <= 1'b0;
            12'h25d: oData <= 1'b0;
            12'h25e: oData <= 1'b0;
            12'h25f: oData <= 1'b0;
            12'h260: oData <= 1'b0;
            12'h261: oData <= 1'b0;
            12'h262: oData <= 1'b0;
            12'h263: oData <= 1'b0;
            12'h264: oData <= 1'b0;
            12'h265: oData <= 1'b0;
            12'h266: oData <= 1'b0;
            12'h267: oData <= 1'b0;
            12'h268: oData <= 1'b0;
            12'h269: oData <= 1'b0;
            12'h26a: oData <= 1'b0;
            12'h26b: oData <= 1'b0;
            12'h26c: oData <= 1'b0;
            12'h26d: oData <= 1'b0;
            12'h26e: oData <= 1'b0;
            12'h26f: oData <= 1'b0;
            12'h270: oData <= 1'b0;
            12'h271: oData <= 1'b0;
            12'h272: oData <= 1'b0;
            12'h273: oData <= 1'b0;
            12'h274: oData <= 1'b0;
            12'h275: oData <= 1'b0;
            12'h276: oData <= 1'b0;
            12'h277: oData <= 1'b0;
            12'h278: oData <= 1'b0;
            12'h279: oData <= 1'b0;
            12'h27a: oData <= 1'b0;
            12'h27b: oData <= 1'b0;
            12'h27c: oData <= 1'b0;
            12'h27d: oData <= 1'b0;
            12'h27e: oData <= 1'b0;
            12'h27f: oData <= 1'b0;
            12'h280: oData <= 1'b0;
            12'h281: oData <= 1'b0;
            12'h282: oData <= 1'b0;
            12'h283: oData <= 1'b0;
            12'h284: oData <= 1'b0;
            12'h285: oData <= 1'b0;
            12'h286: oData <= 1'b0;
            12'h287: oData <= 1'b0;
            12'h288: oData <= 1'b0;
            12'h289: oData <= 1'b0;
            12'h28a: oData <= 1'b0;
            12'h28b: oData <= 1'b0;
            12'h28c: oData <= 1'b0;
            12'h28d: oData <= 1'b0;
            12'h28e: oData <= 1'b0;
            12'h28f: oData <= 1'b0;
            12'h290: oData <= 1'b0;
            12'h291: oData <= 1'b0;
            12'h292: oData <= 1'b0;
            12'h293: oData <= 1'b0;
            12'h294: oData <= 1'b0;
            12'h295: oData <= 1'b0;
            12'h296: oData <= 1'b0;
            12'h297: oData <= 1'b0;
            12'h298: oData <= 1'b0;
            12'h299: oData <= 1'b0;
            12'h29a: oData <= 1'b0;
            12'h29b: oData <= 1'b0;
            12'h29c: oData <= 1'b0;
            12'h29d: oData <= 1'b0;
            12'h29e: oData <= 1'b0;
            12'h29f: oData <= 1'b0;
            12'h2a0: oData <= 1'b0;
            12'h2a1: oData <= 1'b0;
            12'h2a2: oData <= 1'b0;
            12'h2a3: oData <= 1'b0;
            12'h2a4: oData <= 1'b0;
            12'h2a5: oData <= 1'b0;
            12'h2a6: oData <= 1'b0;
            12'h2a7: oData <= 1'b0;
            12'h2a8: oData <= 1'b0;
            12'h2a9: oData <= 1'b0;
            12'h2aa: oData <= 1'b0;
            12'h2ab: oData <= 1'b0;
            12'h2ac: oData <= 1'b0;
            12'h2ad: oData <= 1'b0;
            12'h2ae: oData <= 1'b0;
            12'h2af: oData <= 1'b0;
            12'h2b0: oData <= 1'b0;
            12'h2b1: oData <= 1'b0;
            12'h2b2: oData <= 1'b0;
            12'h2b3: oData <= 1'b0;
            12'h2b4: oData <= 1'b0;
            12'h2b5: oData <= 1'b0;
            12'h2b6: oData <= 1'b0;
            12'h2b7: oData <= 1'b0;
            12'h2b8: oData <= 1'b0;
            12'h2b9: oData <= 1'b0;
            12'h2ba: oData <= 1'b0;
            12'h2bb: oData <= 1'b0;
            12'h2bc: oData <= 1'b0;
            12'h2bd: oData <= 1'b0;
            12'h2be: oData <= 1'b0;
            12'h2bf: oData <= 1'b0;
            12'h2c0: oData <= 1'b0;
            12'h2c1: oData <= 1'b0;
            12'h2c2: oData <= 1'b0;
            12'h2c3: oData <= 1'b0;
            12'h2c4: oData <= 1'b0;
            12'h2c5: oData <= 1'b0;
            12'h2c6: oData <= 1'b0;
            12'h2c7: oData <= 1'b0;
            12'h2c8: oData <= 1'b0;
            12'h2c9: oData <= 1'b0;
            12'h2ca: oData <= 1'b0;
            12'h2cb: oData <= 1'b0;
            12'h2cc: oData <= 1'b0;
            12'h2cd: oData <= 1'b0;
            12'h2ce: oData <= 1'b0;
            12'h2cf: oData <= 1'b0;
            12'h2d0: oData <= 1'b0;
            12'h2d1: oData <= 1'b0;
            12'h2d2: oData <= 1'b0;
            12'h2d3: oData <= 1'b0;
            12'h2d4: oData <= 1'b0;
            12'h2d5: oData <= 1'b0;
            12'h2d6: oData <= 1'b0;
            12'h2d7: oData <= 1'b0;
            12'h2d8: oData <= 1'b0;
            12'h2d9: oData <= 1'b0;
            12'h2da: oData <= 1'b0;
            12'h2db: oData <= 1'b0;
            12'h2dc: oData <= 1'b0;
            12'h2dd: oData <= 1'b0;
            12'h2de: oData <= 1'b0;
            12'h2df: oData <= 1'b0;
            12'h2e0: oData <= 1'b0;
            12'h2e1: oData <= 1'b0;
            12'h2e2: oData <= 1'b0;
            12'h2e3: oData <= 1'b0;
            12'h2e4: oData <= 1'b0;
            12'h2e5: oData <= 1'b0;
            12'h2e6: oData <= 1'b0;
            12'h2e7: oData <= 1'b0;
            12'h2e8: oData <= 1'b0;
            12'h2e9: oData <= 1'b0;
            12'h2ea: oData <= 1'b0;
            12'h2eb: oData <= 1'b0;
            12'h2ec: oData <= 1'b0;
            12'h2ed: oData <= 1'b0;
            12'h2ee: oData <= 1'b0;
            12'h2ef: oData <= 1'b0;
            12'h2f0: oData <= 1'b0;
            12'h2f1: oData <= 1'b0;
            12'h2f2: oData <= 1'b0;
            12'h2f3: oData <= 1'b0;
            12'h2f4: oData <= 1'b0;
            12'h2f5: oData <= 1'b0;
            12'h2f6: oData <= 1'b0;
            12'h2f7: oData <= 1'b0;
            12'h2f8: oData <= 1'b0;
            12'h2f9: oData <= 1'b0;
            12'h2fa: oData <= 1'b0;
            12'h2fb: oData <= 1'b0;
            12'h2fc: oData <= 1'b0;
            12'h2fd: oData <= 1'b0;
            12'h2fe: oData <= 1'b0;
            12'h2ff: oData <= 1'b0;
            12'h300: oData <= 1'b1;
            12'h301: oData <= 1'b1;
            12'h302: oData <= 1'b1;
            12'h303: oData <= 1'b1;
            12'h304: oData <= 1'b0;
            12'h305: oData <= 1'b0;
            12'h306: oData <= 1'b0;
            12'h307: oData <= 1'b0;
            12'h308: oData <= 1'b0;
            12'h309: oData <= 1'b0;
            12'h30a: oData <= 1'b0;
            12'h30b: oData <= 1'b0;
            12'h30c: oData <= 1'b0;
            12'h30d: oData <= 1'b0;
            12'h30e: oData <= 1'b0;
            12'h30f: oData <= 1'b0;
            12'h310: oData <= 1'b1;
            12'h311: oData <= 1'b1;
            12'h312: oData <= 1'b1;
            12'h313: oData <= 1'b1;
            12'h314: oData <= 1'b0;
            12'h315: oData <= 1'b0;
            12'h316: oData <= 1'b0;
            12'h317: oData <= 1'b0;
            12'h318: oData <= 1'b0;
            12'h319: oData <= 1'b0;
            12'h31a: oData <= 1'b0;
            12'h31b: oData <= 1'b0;
            12'h31c: oData <= 1'b0;
            12'h31d: oData <= 1'b0;
            12'h31e: oData <= 1'b0;
            12'h31f: oData <= 1'b0;
            12'h320: oData <= 1'b1;
            12'h321: oData <= 1'b1;
            12'h322: oData <= 1'b1;
            12'h323: oData <= 1'b0;
            12'h324: oData <= 1'b0;
            12'h325: oData <= 1'b0;
            12'h326: oData <= 1'b0;
            12'h327: oData <= 1'b0;
            12'h328: oData <= 1'b0;
            12'h329: oData <= 1'b0;
            12'h32a: oData <= 1'b0;
            12'h32b: oData <= 1'b0;
            12'h32c: oData <= 1'b0;
            12'h32d: oData <= 1'b0;
            12'h32e: oData <= 1'b0;
            12'h32f: oData <= 1'b0;
            12'h330: oData <= 1'b1;
            12'h331: oData <= 1'b1;
            12'h332: oData <= 1'b0;
            12'h333: oData <= 1'b0;
            12'h334: oData <= 1'b0;
            12'h335: oData <= 1'b0;
            12'h336: oData <= 1'b0;
            12'h337: oData <= 1'b0;
            12'h338: oData <= 1'b0;
            12'h339: oData <= 1'b0;
            12'h33a: oData <= 1'b0;
            12'h33b: oData <= 1'b0;
            12'h33c: oData <= 1'b0;
            12'h33d: oData <= 1'b0;
            12'h33e: oData <= 1'b0;
            12'h33f: oData <= 1'b0;
            12'h340: oData <= 1'b0;
            12'h341: oData <= 1'b0;
            12'h342: oData <= 1'b0;
            12'h343: oData <= 1'b0;
            12'h344: oData <= 1'b0;
            12'h345: oData <= 1'b0;
            12'h346: oData <= 1'b0;
            12'h347: oData <= 1'b0;
            12'h348: oData <= 1'b0;
            12'h349: oData <= 1'b0;
            12'h34a: oData <= 1'b0;
            12'h34b: oData <= 1'b0;
            12'h34c: oData <= 1'b0;
            12'h34d: oData <= 1'b0;
            12'h34e: oData <= 1'b0;
            12'h34f: oData <= 1'b0;
            12'h350: oData <= 1'b0;
            12'h351: oData <= 1'b0;
            12'h352: oData <= 1'b0;
            12'h353: oData <= 1'b0;
            12'h354: oData <= 1'b0;
            12'h355: oData <= 1'b0;
            12'h356: oData <= 1'b0;
            12'h357: oData <= 1'b0;
            12'h358: oData <= 1'b0;
            12'h359: oData <= 1'b0;
            12'h35a: oData <= 1'b0;
            12'h35b: oData <= 1'b0;
            12'h35c: oData <= 1'b0;
            12'h35d: oData <= 1'b0;
            12'h35e: oData <= 1'b0;
            12'h35f: oData <= 1'b0;
            12'h360: oData <= 1'b0;
            12'h361: oData <= 1'b0;
            12'h362: oData <= 1'b0;
            12'h363: oData <= 1'b0;
            12'h364: oData <= 1'b0;
            12'h365: oData <= 1'b0;
            12'h366: oData <= 1'b0;
            12'h367: oData <= 1'b0;
            12'h368: oData <= 1'b0;
            12'h369: oData <= 1'b0;
            12'h36a: oData <= 1'b0;
            12'h36b: oData <= 1'b0;
            12'h36c: oData <= 1'b0;
            12'h36d: oData <= 1'b0;
            12'h36e: oData <= 1'b0;
            12'h36f: oData <= 1'b0;
            12'h370: oData <= 1'b0;
            12'h371: oData <= 1'b0;
            12'h372: oData <= 1'b0;
            12'h373: oData <= 1'b0;
            12'h374: oData <= 1'b0;
            12'h375: oData <= 1'b0;
            12'h376: oData <= 1'b0;
            12'h377: oData <= 1'b0;
            12'h378: oData <= 1'b0;
            12'h379: oData <= 1'b0;
            12'h37a: oData <= 1'b0;
            12'h37b: oData <= 1'b0;
            12'h37c: oData <= 1'b0;
            12'h37d: oData <= 1'b0;
            12'h37e: oData <= 1'b0;
            12'h37f: oData <= 1'b0;
            12'h380: oData <= 1'b0;
            12'h381: oData <= 1'b0;
            12'h382: oData <= 1'b0;
            12'h383: oData <= 1'b0;
            12'h384: oData <= 1'b0;
            12'h385: oData <= 1'b0;
            12'h386: oData <= 1'b0;
            12'h387: oData <= 1'b0;
            12'h388: oData <= 1'b0;
            12'h389: oData <= 1'b0;
            12'h38a: oData <= 1'b0;
            12'h38b: oData <= 1'b0;
            12'h38c: oData <= 1'b0;
            12'h38d: oData <= 1'b0;
            12'h38e: oData <= 1'b0;
            12'h38f: oData <= 1'b0;
            12'h390: oData <= 1'b0;
            12'h391: oData <= 1'b0;
            12'h392: oData <= 1'b0;
            12'h393: oData <= 1'b0;
            12'h394: oData <= 1'b0;
            12'h395: oData <= 1'b0;
            12'h396: oData <= 1'b0;
            12'h397: oData <= 1'b0;
            12'h398: oData <= 1'b0;
            12'h399: oData <= 1'b0;
            12'h39a: oData <= 1'b0;
            12'h39b: oData <= 1'b0;
            12'h39c: oData <= 1'b0;
            12'h39d: oData <= 1'b0;
            12'h39e: oData <= 1'b0;
            12'h39f: oData <= 1'b0;
            12'h3a0: oData <= 1'b0;
            12'h3a1: oData <= 1'b0;
            12'h3a2: oData <= 1'b0;
            12'h3a3: oData <= 1'b0;
            12'h3a4: oData <= 1'b0;
            12'h3a5: oData <= 1'b0;
            12'h3a6: oData <= 1'b0;
            12'h3a7: oData <= 1'b0;
            12'h3a8: oData <= 1'b0;
            12'h3a9: oData <= 1'b0;
            12'h3aa: oData <= 1'b0;
            12'h3ab: oData <= 1'b0;
            12'h3ac: oData <= 1'b0;
            12'h3ad: oData <= 1'b0;
            12'h3ae: oData <= 1'b0;
            12'h3af: oData <= 1'b0;
            12'h3b0: oData <= 1'b0;
            12'h3b1: oData <= 1'b0;
            12'h3b2: oData <= 1'b0;
            12'h3b3: oData <= 1'b0;
            12'h3b4: oData <= 1'b0;
            12'h3b5: oData <= 1'b0;
            12'h3b6: oData <= 1'b0;
            12'h3b7: oData <= 1'b0;
            12'h3b8: oData <= 1'b0;
            12'h3b9: oData <= 1'b0;
            12'h3ba: oData <= 1'b0;
            12'h3bb: oData <= 1'b0;
            12'h3bc: oData <= 1'b0;
            12'h3bd: oData <= 1'b0;
            12'h3be: oData <= 1'b0;
            12'h3bf: oData <= 1'b0;
            12'h3c0: oData <= 1'b0;
            12'h3c1: oData <= 1'b0;
            12'h3c2: oData <= 1'b0;
            12'h3c3: oData <= 1'b0;
            12'h3c4: oData <= 1'b0;
            12'h3c5: oData <= 1'b0;
            12'h3c6: oData <= 1'b0;
            12'h3c7: oData <= 1'b0;
            12'h3c8: oData <= 1'b0;
            12'h3c9: oData <= 1'b0;
            12'h3ca: oData <= 1'b0;
            12'h3cb: oData <= 1'b0;
            12'h3cc: oData <= 1'b0;
            12'h3cd: oData <= 1'b0;
            12'h3ce: oData <= 1'b0;
            12'h3cf: oData <= 1'b0;
            12'h3d0: oData <= 1'b0;
            12'h3d1: oData <= 1'b0;
            12'h3d2: oData <= 1'b0;
            12'h3d3: oData <= 1'b0;
            12'h3d4: oData <= 1'b0;
            12'h3d5: oData <= 1'b0;
            12'h3d6: oData <= 1'b0;
            12'h3d7: oData <= 1'b0;
            12'h3d8: oData <= 1'b0;
            12'h3d9: oData <= 1'b0;
            12'h3da: oData <= 1'b0;
            12'h3db: oData <= 1'b0;
            12'h3dc: oData <= 1'b0;
            12'h3dd: oData <= 1'b0;
            12'h3de: oData <= 1'b0;
            12'h3df: oData <= 1'b0;
            12'h3e0: oData <= 1'b0;
            12'h3e1: oData <= 1'b0;
            12'h3e2: oData <= 1'b0;
            12'h3e3: oData <= 1'b0;
            12'h3e4: oData <= 1'b0;
            12'h3e5: oData <= 1'b0;
            12'h3e6: oData <= 1'b0;
            12'h3e7: oData <= 1'b0;
            12'h3e8: oData <= 1'b0;
            12'h3e9: oData <= 1'b0;
            12'h3ea: oData <= 1'b0;
            12'h3eb: oData <= 1'b0;
            12'h3ec: oData <= 1'b0;
            12'h3ed: oData <= 1'b0;
            12'h3ee: oData <= 1'b0;
            12'h3ef: oData <= 1'b0;
            12'h3f0: oData <= 1'b0;
            12'h3f1: oData <= 1'b0;
            12'h3f2: oData <= 1'b0;
            12'h3f3: oData <= 1'b0;
            12'h3f4: oData <= 1'b0;
            12'h3f5: oData <= 1'b0;
            12'h3f6: oData <= 1'b0;
            12'h3f7: oData <= 1'b0;
            12'h3f8: oData <= 1'b0;
            12'h3f9: oData <= 1'b0;
            12'h3fa: oData <= 1'b0;
            12'h3fb: oData <= 1'b0;
            12'h3fc: oData <= 1'b0;
            12'h3fd: oData <= 1'b0;
            12'h3fe: oData <= 1'b0;
            12'h3ff: oData <= 1'b0;
            12'h400: oData <= 1'b1;
            12'h401: oData <= 1'b1;
            12'h402: oData <= 1'b1;
            12'h403: oData <= 1'b1;
            12'h404: oData <= 1'b1;
            12'h405: oData <= 1'b0;
            12'h406: oData <= 1'b0;
            12'h407: oData <= 1'b0;
            12'h408: oData <= 1'b0;
            12'h409: oData <= 1'b0;
            12'h40a: oData <= 1'b0;
            12'h40b: oData <= 1'b0;
            12'h40c: oData <= 1'b0;
            12'h40d: oData <= 1'b0;
            12'h40e: oData <= 1'b0;
            12'h40f: oData <= 1'b0;
            12'h410: oData <= 1'b1;
            12'h411: oData <= 1'b1;
            12'h412: oData <= 1'b1;
            12'h413: oData <= 1'b1;
            12'h414: oData <= 1'b1;
            12'h415: oData <= 1'b0;
            12'h416: oData <= 1'b0;
            12'h417: oData <= 1'b0;
            12'h418: oData <= 1'b0;
            12'h419: oData <= 1'b0;
            12'h41a: oData <= 1'b0;
            12'h41b: oData <= 1'b0;
            12'h41c: oData <= 1'b0;
            12'h41d: oData <= 1'b0;
            12'h41e: oData <= 1'b0;
            12'h41f: oData <= 1'b0;
            12'h420: oData <= 1'b1;
            12'h421: oData <= 1'b1;
            12'h422: oData <= 1'b1;
            12'h423: oData <= 1'b1;
            12'h424: oData <= 1'b0;
            12'h425: oData <= 1'b0;
            12'h426: oData <= 1'b0;
            12'h427: oData <= 1'b0;
            12'h428: oData <= 1'b0;
            12'h429: oData <= 1'b0;
            12'h42a: oData <= 1'b0;
            12'h42b: oData <= 1'b0;
            12'h42c: oData <= 1'b0;
            12'h42d: oData <= 1'b0;
            12'h42e: oData <= 1'b0;
            12'h42f: oData <= 1'b0;
            12'h430: oData <= 1'b1;
            12'h431: oData <= 1'b1;
            12'h432: oData <= 1'b1;
            12'h433: oData <= 1'b0;
            12'h434: oData <= 1'b0;
            12'h435: oData <= 1'b0;
            12'h436: oData <= 1'b0;
            12'h437: oData <= 1'b0;
            12'h438: oData <= 1'b0;
            12'h439: oData <= 1'b0;
            12'h43a: oData <= 1'b0;
            12'h43b: oData <= 1'b0;
            12'h43c: oData <= 1'b0;
            12'h43d: oData <= 1'b0;
            12'h43e: oData <= 1'b0;
            12'h43f: oData <= 1'b0;
            12'h440: oData <= 1'b1;
            12'h441: oData <= 1'b1;
            12'h442: oData <= 1'b0;
            12'h443: oData <= 1'b0;
            12'h444: oData <= 1'b0;
            12'h445: oData <= 1'b0;
            12'h446: oData <= 1'b0;
            12'h447: oData <= 1'b0;
            12'h448: oData <= 1'b0;
            12'h449: oData <= 1'b0;
            12'h44a: oData <= 1'b0;
            12'h44b: oData <= 1'b0;
            12'h44c: oData <= 1'b0;
            12'h44d: oData <= 1'b0;
            12'h44e: oData <= 1'b0;
            12'h44f: oData <= 1'b0;
            12'h450: oData <= 1'b0;
            12'h451: oData <= 1'b0;
            12'h452: oData <= 1'b0;
            12'h453: oData <= 1'b0;
            12'h454: oData <= 1'b0;
            12'h455: oData <= 1'b0;
            12'h456: oData <= 1'b0;
            12'h457: oData <= 1'b0;
            12'h458: oData <= 1'b0;
            12'h459: oData <= 1'b0;
            12'h45a: oData <= 1'b0;
            12'h45b: oData <= 1'b0;
            12'h45c: oData <= 1'b0;
            12'h45d: oData <= 1'b0;
            12'h45e: oData <= 1'b0;
            12'h45f: oData <= 1'b0;
            12'h460: oData <= 1'b0;
            12'h461: oData <= 1'b0;
            12'h462: oData <= 1'b0;
            12'h463: oData <= 1'b0;
            12'h464: oData <= 1'b0;
            12'h465: oData <= 1'b0;
            12'h466: oData <= 1'b0;
            12'h467: oData <= 1'b0;
            12'h468: oData <= 1'b0;
            12'h469: oData <= 1'b0;
            12'h46a: oData <= 1'b0;
            12'h46b: oData <= 1'b0;
            12'h46c: oData <= 1'b0;
            12'h46d: oData <= 1'b0;
            12'h46e: oData <= 1'b0;
            12'h46f: oData <= 1'b0;
            12'h470: oData <= 1'b0;
            12'h471: oData <= 1'b0;
            12'h472: oData <= 1'b0;
            12'h473: oData <= 1'b0;
            12'h474: oData <= 1'b0;
            12'h475: oData <= 1'b0;
            12'h476: oData <= 1'b0;
            12'h477: oData <= 1'b0;
            12'h478: oData <= 1'b0;
            12'h479: oData <= 1'b0;
            12'h47a: oData <= 1'b0;
            12'h47b: oData <= 1'b0;
            12'h47c: oData <= 1'b0;
            12'h47d: oData <= 1'b0;
            12'h47e: oData <= 1'b0;
            12'h47f: oData <= 1'b0;
            12'h480: oData <= 1'b0;
            12'h481: oData <= 1'b0;
            12'h482: oData <= 1'b0;
            12'h483: oData <= 1'b0;
            12'h484: oData <= 1'b0;
            12'h485: oData <= 1'b0;
            12'h486: oData <= 1'b0;
            12'h487: oData <= 1'b0;
            12'h488: oData <= 1'b0;
            12'h489: oData <= 1'b0;
            12'h48a: oData <= 1'b0;
            12'h48b: oData <= 1'b0;
            12'h48c: oData <= 1'b0;
            12'h48d: oData <= 1'b0;
            12'h48e: oData <= 1'b0;
            12'h48f: oData <= 1'b0;
            12'h490: oData <= 1'b0;
            12'h491: oData <= 1'b0;
            12'h492: oData <= 1'b0;
            12'h493: oData <= 1'b0;
            12'h494: oData <= 1'b0;
            12'h495: oData <= 1'b0;
            12'h496: oData <= 1'b0;
            12'h497: oData <= 1'b0;
            12'h498: oData <= 1'b0;
            12'h499: oData <= 1'b0;
            12'h49a: oData <= 1'b0;
            12'h49b: oData <= 1'b0;
            12'h49c: oData <= 1'b0;
            12'h49d: oData <= 1'b0;
            12'h49e: oData <= 1'b0;
            12'h49f: oData <= 1'b0;
            12'h4a0: oData <= 1'b0;
            12'h4a1: oData <= 1'b0;
            12'h4a2: oData <= 1'b0;
            12'h4a3: oData <= 1'b0;
            12'h4a4: oData <= 1'b0;
            12'h4a5: oData <= 1'b0;
            12'h4a6: oData <= 1'b0;
            12'h4a7: oData <= 1'b0;
            12'h4a8: oData <= 1'b0;
            12'h4a9: oData <= 1'b0;
            12'h4aa: oData <= 1'b0;
            12'h4ab: oData <= 1'b0;
            12'h4ac: oData <= 1'b0;
            12'h4ad: oData <= 1'b0;
            12'h4ae: oData <= 1'b0;
            12'h4af: oData <= 1'b0;
            12'h4b0: oData <= 1'b0;
            12'h4b1: oData <= 1'b0;
            12'h4b2: oData <= 1'b0;
            12'h4b3: oData <= 1'b0;
            12'h4b4: oData <= 1'b0;
            12'h4b5: oData <= 1'b0;
            12'h4b6: oData <= 1'b0;
            12'h4b7: oData <= 1'b0;
            12'h4b8: oData <= 1'b0;
            12'h4b9: oData <= 1'b0;
            12'h4ba: oData <= 1'b0;
            12'h4bb: oData <= 1'b0;
            12'h4bc: oData <= 1'b0;
            12'h4bd: oData <= 1'b0;
            12'h4be: oData <= 1'b0;
            12'h4bf: oData <= 1'b0;
            12'h4c0: oData <= 1'b0;
            12'h4c1: oData <= 1'b0;
            12'h4c2: oData <= 1'b0;
            12'h4c3: oData <= 1'b0;
            12'h4c4: oData <= 1'b0;
            12'h4c5: oData <= 1'b0;
            12'h4c6: oData <= 1'b0;
            12'h4c7: oData <= 1'b0;
            12'h4c8: oData <= 1'b0;
            12'h4c9: oData <= 1'b0;
            12'h4ca: oData <= 1'b0;
            12'h4cb: oData <= 1'b0;
            12'h4cc: oData <= 1'b0;
            12'h4cd: oData <= 1'b0;
            12'h4ce: oData <= 1'b0;
            12'h4cf: oData <= 1'b0;
            12'h4d0: oData <= 1'b0;
            12'h4d1: oData <= 1'b0;
            12'h4d2: oData <= 1'b0;
            12'h4d3: oData <= 1'b0;
            12'h4d4: oData <= 1'b0;
            12'h4d5: oData <= 1'b0;
            12'h4d6: oData <= 1'b0;
            12'h4d7: oData <= 1'b0;
            12'h4d8: oData <= 1'b0;
            12'h4d9: oData <= 1'b0;
            12'h4da: oData <= 1'b0;
            12'h4db: oData <= 1'b0;
            12'h4dc: oData <= 1'b0;
            12'h4dd: oData <= 1'b0;
            12'h4de: oData <= 1'b0;
            12'h4df: oData <= 1'b0;
            12'h4e0: oData <= 1'b0;
            12'h4e1: oData <= 1'b0;
            12'h4e2: oData <= 1'b0;
            12'h4e3: oData <= 1'b0;
            12'h4e4: oData <= 1'b0;
            12'h4e5: oData <= 1'b0;
            12'h4e6: oData <= 1'b0;
            12'h4e7: oData <= 1'b0;
            12'h4e8: oData <= 1'b0;
            12'h4e9: oData <= 1'b0;
            12'h4ea: oData <= 1'b0;
            12'h4eb: oData <= 1'b0;
            12'h4ec: oData <= 1'b0;
            12'h4ed: oData <= 1'b0;
            12'h4ee: oData <= 1'b0;
            12'h4ef: oData <= 1'b0;
            12'h4f0: oData <= 1'b0;
            12'h4f1: oData <= 1'b0;
            12'h4f2: oData <= 1'b0;
            12'h4f3: oData <= 1'b0;
            12'h4f4: oData <= 1'b0;
            12'h4f5: oData <= 1'b0;
            12'h4f6: oData <= 1'b0;
            12'h4f7: oData <= 1'b0;
            12'h4f8: oData <= 1'b0;
            12'h4f9: oData <= 1'b0;
            12'h4fa: oData <= 1'b0;
            12'h4fb: oData <= 1'b0;
            12'h4fc: oData <= 1'b0;
            12'h4fd: oData <= 1'b0;
            12'h4fe: oData <= 1'b0;
            12'h4ff: oData <= 1'b0;
            12'h500: oData <= 1'b1;
            12'h501: oData <= 1'b1;
            12'h502: oData <= 1'b1;
            12'h503: oData <= 1'b1;
            12'h504: oData <= 1'b1;
            12'h505: oData <= 1'b1;
            12'h506: oData <= 1'b0;
            12'h507: oData <= 1'b0;
            12'h508: oData <= 1'b0;
            12'h509: oData <= 1'b0;
            12'h50a: oData <= 1'b0;
            12'h50b: oData <= 1'b0;
            12'h50c: oData <= 1'b0;
            12'h50d: oData <= 1'b0;
            12'h50e: oData <= 1'b0;
            12'h50f: oData <= 1'b0;
            12'h510: oData <= 1'b1;
            12'h511: oData <= 1'b1;
            12'h512: oData <= 1'b1;
            12'h513: oData <= 1'b1;
            12'h514: oData <= 1'b1;
            12'h515: oData <= 1'b1;
            12'h516: oData <= 1'b0;
            12'h517: oData <= 1'b0;
            12'h518: oData <= 1'b0;
            12'h519: oData <= 1'b0;
            12'h51a: oData <= 1'b0;
            12'h51b: oData <= 1'b0;
            12'h51c: oData <= 1'b0;
            12'h51d: oData <= 1'b0;
            12'h51e: oData <= 1'b0;
            12'h51f: oData <= 1'b0;
            12'h520: oData <= 1'b1;
            12'h521: oData <= 1'b1;
            12'h522: oData <= 1'b1;
            12'h523: oData <= 1'b1;
            12'h524: oData <= 1'b1;
            12'h525: oData <= 1'b0;
            12'h526: oData <= 1'b0;
            12'h527: oData <= 1'b0;
            12'h528: oData <= 1'b0;
            12'h529: oData <= 1'b0;
            12'h52a: oData <= 1'b0;
            12'h52b: oData <= 1'b0;
            12'h52c: oData <= 1'b0;
            12'h52d: oData <= 1'b0;
            12'h52e: oData <= 1'b0;
            12'h52f: oData <= 1'b0;
            12'h530: oData <= 1'b1;
            12'h531: oData <= 1'b1;
            12'h532: oData <= 1'b1;
            12'h533: oData <= 1'b1;
            12'h534: oData <= 1'b1;
            12'h535: oData <= 1'b0;
            12'h536: oData <= 1'b0;
            12'h537: oData <= 1'b0;
            12'h538: oData <= 1'b0;
            12'h539: oData <= 1'b0;
            12'h53a: oData <= 1'b0;
            12'h53b: oData <= 1'b0;
            12'h53c: oData <= 1'b0;
            12'h53d: oData <= 1'b0;
            12'h53e: oData <= 1'b0;
            12'h53f: oData <= 1'b0;
            12'h540: oData <= 1'b1;
            12'h541: oData <= 1'b1;
            12'h542: oData <= 1'b1;
            12'h543: oData <= 1'b1;
            12'h544: oData <= 1'b0;
            12'h545: oData <= 1'b0;
            12'h546: oData <= 1'b0;
            12'h547: oData <= 1'b0;
            12'h548: oData <= 1'b0;
            12'h549: oData <= 1'b0;
            12'h54a: oData <= 1'b0;
            12'h54b: oData <= 1'b0;
            12'h54c: oData <= 1'b0;
            12'h54d: oData <= 1'b0;
            12'h54e: oData <= 1'b0;
            12'h54f: oData <= 1'b0;
            12'h550: oData <= 1'b1;
            12'h551: oData <= 1'b1;
            12'h552: oData <= 1'b0;
            12'h553: oData <= 1'b0;
            12'h554: oData <= 1'b0;
            12'h555: oData <= 1'b0;
            12'h556: oData <= 1'b0;
            12'h557: oData <= 1'b0;
            12'h558: oData <= 1'b0;
            12'h559: oData <= 1'b0;
            12'h55a: oData <= 1'b0;
            12'h55b: oData <= 1'b0;
            12'h55c: oData <= 1'b0;
            12'h55d: oData <= 1'b0;
            12'h55e: oData <= 1'b0;
            12'h55f: oData <= 1'b0;
            12'h560: oData <= 1'b0;
            12'h561: oData <= 1'b0;
            12'h562: oData <= 1'b0;
            12'h563: oData <= 1'b0;
            12'h564: oData <= 1'b0;
            12'h565: oData <= 1'b0;
            12'h566: oData <= 1'b0;
            12'h567: oData <= 1'b0;
            12'h568: oData <= 1'b0;
            12'h569: oData <= 1'b0;
            12'h56a: oData <= 1'b0;
            12'h56b: oData <= 1'b0;
            12'h56c: oData <= 1'b0;
            12'h56d: oData <= 1'b0;
            12'h56e: oData <= 1'b0;
            12'h56f: oData <= 1'b0;
            12'h570: oData <= 1'b0;
            12'h571: oData <= 1'b0;
            12'h572: oData <= 1'b0;
            12'h573: oData <= 1'b0;
            12'h574: oData <= 1'b0;
            12'h575: oData <= 1'b0;
            12'h576: oData <= 1'b0;
            12'h577: oData <= 1'b0;
            12'h578: oData <= 1'b0;
            12'h579: oData <= 1'b0;
            12'h57a: oData <= 1'b0;
            12'h57b: oData <= 1'b0;
            12'h57c: oData <= 1'b0;
            12'h57d: oData <= 1'b0;
            12'h57e: oData <= 1'b0;
            12'h57f: oData <= 1'b0;
            12'h580: oData <= 1'b0;
            12'h581: oData <= 1'b0;
            12'h582: oData <= 1'b0;
            12'h583: oData <= 1'b0;
            12'h584: oData <= 1'b0;
            12'h585: oData <= 1'b0;
            12'h586: oData <= 1'b0;
            12'h587: oData <= 1'b0;
            12'h588: oData <= 1'b0;
            12'h589: oData <= 1'b0;
            12'h58a: oData <= 1'b0;
            12'h58b: oData <= 1'b0;
            12'h58c: oData <= 1'b0;
            12'h58d: oData <= 1'b0;
            12'h58e: oData <= 1'b0;
            12'h58f: oData <= 1'b0;
            12'h590: oData <= 1'b0;
            12'h591: oData <= 1'b0;
            12'h592: oData <= 1'b0;
            12'h593: oData <= 1'b0;
            12'h594: oData <= 1'b0;
            12'h595: oData <= 1'b0;
            12'h596: oData <= 1'b0;
            12'h597: oData <= 1'b0;
            12'h598: oData <= 1'b0;
            12'h599: oData <= 1'b0;
            12'h59a: oData <= 1'b0;
            12'h59b: oData <= 1'b0;
            12'h59c: oData <= 1'b0;
            12'h59d: oData <= 1'b0;
            12'h59e: oData <= 1'b0;
            12'h59f: oData <= 1'b0;
            12'h5a0: oData <= 1'b0;
            12'h5a1: oData <= 1'b0;
            12'h5a2: oData <= 1'b0;
            12'h5a3: oData <= 1'b0;
            12'h5a4: oData <= 1'b0;
            12'h5a5: oData <= 1'b0;
            12'h5a6: oData <= 1'b0;
            12'h5a7: oData <= 1'b0;
            12'h5a8: oData <= 1'b0;
            12'h5a9: oData <= 1'b0;
            12'h5aa: oData <= 1'b0;
            12'h5ab: oData <= 1'b0;
            12'h5ac: oData <= 1'b0;
            12'h5ad: oData <= 1'b0;
            12'h5ae: oData <= 1'b0;
            12'h5af: oData <= 1'b0;
            12'h5b0: oData <= 1'b0;
            12'h5b1: oData <= 1'b0;
            12'h5b2: oData <= 1'b0;
            12'h5b3: oData <= 1'b0;
            12'h5b4: oData <= 1'b0;
            12'h5b5: oData <= 1'b0;
            12'h5b6: oData <= 1'b0;
            12'h5b7: oData <= 1'b0;
            12'h5b8: oData <= 1'b0;
            12'h5b9: oData <= 1'b0;
            12'h5ba: oData <= 1'b0;
            12'h5bb: oData <= 1'b0;
            12'h5bc: oData <= 1'b0;
            12'h5bd: oData <= 1'b0;
            12'h5be: oData <= 1'b0;
            12'h5bf: oData <= 1'b0;
            12'h5c0: oData <= 1'b0;
            12'h5c1: oData <= 1'b0;
            12'h5c2: oData <= 1'b0;
            12'h5c3: oData <= 1'b0;
            12'h5c4: oData <= 1'b0;
            12'h5c5: oData <= 1'b0;
            12'h5c6: oData <= 1'b0;
            12'h5c7: oData <= 1'b0;
            12'h5c8: oData <= 1'b0;
            12'h5c9: oData <= 1'b0;
            12'h5ca: oData <= 1'b0;
            12'h5cb: oData <= 1'b0;
            12'h5cc: oData <= 1'b0;
            12'h5cd: oData <= 1'b0;
            12'h5ce: oData <= 1'b0;
            12'h5cf: oData <= 1'b0;
            12'h5d0: oData <= 1'b0;
            12'h5d1: oData <= 1'b0;
            12'h5d2: oData <= 1'b0;
            12'h5d3: oData <= 1'b0;
            12'h5d4: oData <= 1'b0;
            12'h5d5: oData <= 1'b0;
            12'h5d6: oData <= 1'b0;
            12'h5d7: oData <= 1'b0;
            12'h5d8: oData <= 1'b0;
            12'h5d9: oData <= 1'b0;
            12'h5da: oData <= 1'b0;
            12'h5db: oData <= 1'b0;
            12'h5dc: oData <= 1'b0;
            12'h5dd: oData <= 1'b0;
            12'h5de: oData <= 1'b0;
            12'h5df: oData <= 1'b0;
            12'h5e0: oData <= 1'b0;
            12'h5e1: oData <= 1'b0;
            12'h5e2: oData <= 1'b0;
            12'h5e3: oData <= 1'b0;
            12'h5e4: oData <= 1'b0;
            12'h5e5: oData <= 1'b0;
            12'h5e6: oData <= 1'b0;
            12'h5e7: oData <= 1'b0;
            12'h5e8: oData <= 1'b0;
            12'h5e9: oData <= 1'b0;
            12'h5ea: oData <= 1'b0;
            12'h5eb: oData <= 1'b0;
            12'h5ec: oData <= 1'b0;
            12'h5ed: oData <= 1'b0;
            12'h5ee: oData <= 1'b0;
            12'h5ef: oData <= 1'b0;
            12'h5f0: oData <= 1'b0;
            12'h5f1: oData <= 1'b0;
            12'h5f2: oData <= 1'b0;
            12'h5f3: oData <= 1'b0;
            12'h5f4: oData <= 1'b0;
            12'h5f5: oData <= 1'b0;
            12'h5f6: oData <= 1'b0;
            12'h5f7: oData <= 1'b0;
            12'h5f8: oData <= 1'b0;
            12'h5f9: oData <= 1'b0;
            12'h5fa: oData <= 1'b0;
            12'h5fb: oData <= 1'b0;
            12'h5fc: oData <= 1'b0;
            12'h5fd: oData <= 1'b0;
            12'h5fe: oData <= 1'b0;
            12'h5ff: oData <= 1'b0;
            12'h600: oData <= 1'b1;
            12'h601: oData <= 1'b1;
            12'h602: oData <= 1'b1;
            12'h603: oData <= 1'b1;
            12'h604: oData <= 1'b1;
            12'h605: oData <= 1'b1;
            12'h606: oData <= 1'b1;
            12'h607: oData <= 1'b0;
            12'h608: oData <= 1'b0;
            12'h609: oData <= 1'b0;
            12'h60a: oData <= 1'b0;
            12'h60b: oData <= 1'b0;
            12'h60c: oData <= 1'b0;
            12'h60d: oData <= 1'b0;
            12'h60e: oData <= 1'b0;
            12'h60f: oData <= 1'b0;
            12'h610: oData <= 1'b1;
            12'h611: oData <= 1'b1;
            12'h612: oData <= 1'b1;
            12'h613: oData <= 1'b1;
            12'h614: oData <= 1'b1;
            12'h615: oData <= 1'b1;
            12'h616: oData <= 1'b1;
            12'h617: oData <= 1'b0;
            12'h618: oData <= 1'b0;
            12'h619: oData <= 1'b0;
            12'h61a: oData <= 1'b0;
            12'h61b: oData <= 1'b0;
            12'h61c: oData <= 1'b0;
            12'h61d: oData <= 1'b0;
            12'h61e: oData <= 1'b0;
            12'h61f: oData <= 1'b0;
            12'h620: oData <= 1'b1;
            12'h621: oData <= 1'b1;
            12'h622: oData <= 1'b1;
            12'h623: oData <= 1'b1;
            12'h624: oData <= 1'b1;
            12'h625: oData <= 1'b1;
            12'h626: oData <= 1'b0;
            12'h627: oData <= 1'b0;
            12'h628: oData <= 1'b0;
            12'h629: oData <= 1'b0;
            12'h62a: oData <= 1'b0;
            12'h62b: oData <= 1'b0;
            12'h62c: oData <= 1'b0;
            12'h62d: oData <= 1'b0;
            12'h62e: oData <= 1'b0;
            12'h62f: oData <= 1'b0;
            12'h630: oData <= 1'b1;
            12'h631: oData <= 1'b1;
            12'h632: oData <= 1'b1;
            12'h633: oData <= 1'b1;
            12'h634: oData <= 1'b1;
            12'h635: oData <= 1'b1;
            12'h636: oData <= 1'b0;
            12'h637: oData <= 1'b0;
            12'h638: oData <= 1'b0;
            12'h639: oData <= 1'b0;
            12'h63a: oData <= 1'b0;
            12'h63b: oData <= 1'b0;
            12'h63c: oData <= 1'b0;
            12'h63d: oData <= 1'b0;
            12'h63e: oData <= 1'b0;
            12'h63f: oData <= 1'b0;
            12'h640: oData <= 1'b1;
            12'h641: oData <= 1'b1;
            12'h642: oData <= 1'b1;
            12'h643: oData <= 1'b1;
            12'h644: oData <= 1'b1;
            12'h645: oData <= 1'b0;
            12'h646: oData <= 1'b0;
            12'h647: oData <= 1'b0;
            12'h648: oData <= 1'b0;
            12'h649: oData <= 1'b0;
            12'h64a: oData <= 1'b0;
            12'h64b: oData <= 1'b0;
            12'h64c: oData <= 1'b0;
            12'h64d: oData <= 1'b0;
            12'h64e: oData <= 1'b0;
            12'h64f: oData <= 1'b0;
            12'h650: oData <= 1'b1;
            12'h651: oData <= 1'b1;
            12'h652: oData <= 1'b1;
            12'h653: oData <= 1'b1;
            12'h654: oData <= 1'b0;
            12'h655: oData <= 1'b0;
            12'h656: oData <= 1'b0;
            12'h657: oData <= 1'b0;
            12'h658: oData <= 1'b0;
            12'h659: oData <= 1'b0;
            12'h65a: oData <= 1'b0;
            12'h65b: oData <= 1'b0;
            12'h65c: oData <= 1'b0;
            12'h65d: oData <= 1'b0;
            12'h65e: oData <= 1'b0;
            12'h65f: oData <= 1'b0;
            12'h660: oData <= 1'b1;
            12'h661: oData <= 1'b1;
            12'h662: oData <= 1'b0;
            12'h663: oData <= 1'b0;
            12'h664: oData <= 1'b0;
            12'h665: oData <= 1'b0;
            12'h666: oData <= 1'b0;
            12'h667: oData <= 1'b0;
            12'h668: oData <= 1'b0;
            12'h669: oData <= 1'b0;
            12'h66a: oData <= 1'b0;
            12'h66b: oData <= 1'b0;
            12'h66c: oData <= 1'b0;
            12'h66d: oData <= 1'b0;
            12'h66e: oData <= 1'b0;
            12'h66f: oData <= 1'b0;
            12'h670: oData <= 1'b0;
            12'h671: oData <= 1'b0;
            12'h672: oData <= 1'b0;
            12'h673: oData <= 1'b0;
            12'h674: oData <= 1'b0;
            12'h675: oData <= 1'b0;
            12'h676: oData <= 1'b0;
            12'h677: oData <= 1'b0;
            12'h678: oData <= 1'b0;
            12'h679: oData <= 1'b0;
            12'h67a: oData <= 1'b0;
            12'h67b: oData <= 1'b0;
            12'h67c: oData <= 1'b0;
            12'h67d: oData <= 1'b0;
            12'h67e: oData <= 1'b0;
            12'h67f: oData <= 1'b0;
            12'h680: oData <= 1'b0;
            12'h681: oData <= 1'b0;
            12'h682: oData <= 1'b0;
            12'h683: oData <= 1'b0;
            12'h684: oData <= 1'b0;
            12'h685: oData <= 1'b0;
            12'h686: oData <= 1'b0;
            12'h687: oData <= 1'b0;
            12'h688: oData <= 1'b0;
            12'h689: oData <= 1'b0;
            12'h68a: oData <= 1'b0;
            12'h68b: oData <= 1'b0;
            12'h68c: oData <= 1'b0;
            12'h68d: oData <= 1'b0;
            12'h68e: oData <= 1'b0;
            12'h68f: oData <= 1'b0;
            12'h690: oData <= 1'b0;
            12'h691: oData <= 1'b0;
            12'h692: oData <= 1'b0;
            12'h693: oData <= 1'b0;
            12'h694: oData <= 1'b0;
            12'h695: oData <= 1'b0;
            12'h696: oData <= 1'b0;
            12'h697: oData <= 1'b0;
            12'h698: oData <= 1'b0;
            12'h699: oData <= 1'b0;
            12'h69a: oData <= 1'b0;
            12'h69b: oData <= 1'b0;
            12'h69c: oData <= 1'b0;
            12'h69d: oData <= 1'b0;
            12'h69e: oData <= 1'b0;
            12'h69f: oData <= 1'b0;
            12'h6a0: oData <= 1'b0;
            12'h6a1: oData <= 1'b0;
            12'h6a2: oData <= 1'b0;
            12'h6a3: oData <= 1'b0;
            12'h6a4: oData <= 1'b0;
            12'h6a5: oData <= 1'b0;
            12'h6a6: oData <= 1'b0;
            12'h6a7: oData <= 1'b0;
            12'h6a8: oData <= 1'b0;
            12'h6a9: oData <= 1'b0;
            12'h6aa: oData <= 1'b0;
            12'h6ab: oData <= 1'b0;
            12'h6ac: oData <= 1'b0;
            12'h6ad: oData <= 1'b0;
            12'h6ae: oData <= 1'b0;
            12'h6af: oData <= 1'b0;
            12'h6b0: oData <= 1'b0;
            12'h6b1: oData <= 1'b0;
            12'h6b2: oData <= 1'b0;
            12'h6b3: oData <= 1'b0;
            12'h6b4: oData <= 1'b0;
            12'h6b5: oData <= 1'b0;
            12'h6b6: oData <= 1'b0;
            12'h6b7: oData <= 1'b0;
            12'h6b8: oData <= 1'b0;
            12'h6b9: oData <= 1'b0;
            12'h6ba: oData <= 1'b0;
            12'h6bb: oData <= 1'b0;
            12'h6bc: oData <= 1'b0;
            12'h6bd: oData <= 1'b0;
            12'h6be: oData <= 1'b0;
            12'h6bf: oData <= 1'b0;
            12'h6c0: oData <= 1'b0;
            12'h6c1: oData <= 1'b0;
            12'h6c2: oData <= 1'b0;
            12'h6c3: oData <= 1'b0;
            12'h6c4: oData <= 1'b0;
            12'h6c5: oData <= 1'b0;
            12'h6c6: oData <= 1'b0;
            12'h6c7: oData <= 1'b0;
            12'h6c8: oData <= 1'b0;
            12'h6c9: oData <= 1'b0;
            12'h6ca: oData <= 1'b0;
            12'h6cb: oData <= 1'b0;
            12'h6cc: oData <= 1'b0;
            12'h6cd: oData <= 1'b0;
            12'h6ce: oData <= 1'b0;
            12'h6cf: oData <= 1'b0;
            12'h6d0: oData <= 1'b0;
            12'h6d1: oData <= 1'b0;
            12'h6d2: oData <= 1'b0;
            12'h6d3: oData <= 1'b0;
            12'h6d4: oData <= 1'b0;
            12'h6d5: oData <= 1'b0;
            12'h6d6: oData <= 1'b0;
            12'h6d7: oData <= 1'b0;
            12'h6d8: oData <= 1'b0;
            12'h6d9: oData <= 1'b0;
            12'h6da: oData <= 1'b0;
            12'h6db: oData <= 1'b0;
            12'h6dc: oData <= 1'b0;
            12'h6dd: oData <= 1'b0;
            12'h6de: oData <= 1'b0;
            12'h6df: oData <= 1'b0;
            12'h6e0: oData <= 1'b0;
            12'h6e1: oData <= 1'b0;
            12'h6e2: oData <= 1'b0;
            12'h6e3: oData <= 1'b0;
            12'h6e4: oData <= 1'b0;
            12'h6e5: oData <= 1'b0;
            12'h6e6: oData <= 1'b0;
            12'h6e7: oData <= 1'b0;
            12'h6e8: oData <= 1'b0;
            12'h6e9: oData <= 1'b0;
            12'h6ea: oData <= 1'b0;
            12'h6eb: oData <= 1'b0;
            12'h6ec: oData <= 1'b0;
            12'h6ed: oData <= 1'b0;
            12'h6ee: oData <= 1'b0;
            12'h6ef: oData <= 1'b0;
            12'h6f0: oData <= 1'b0;
            12'h6f1: oData <= 1'b0;
            12'h6f2: oData <= 1'b0;
            12'h6f3: oData <= 1'b0;
            12'h6f4: oData <= 1'b0;
            12'h6f5: oData <= 1'b0;
            12'h6f6: oData <= 1'b0;
            12'h6f7: oData <= 1'b0;
            12'h6f8: oData <= 1'b0;
            12'h6f9: oData <= 1'b0;
            12'h6fa: oData <= 1'b0;
            12'h6fb: oData <= 1'b0;
            12'h6fc: oData <= 1'b0;
            12'h6fd: oData <= 1'b0;
            12'h6fe: oData <= 1'b0;
            12'h6ff: oData <= 1'b0;
            12'h700: oData <= 1'b1;
            12'h701: oData <= 1'b1;
            12'h702: oData <= 1'b1;
            12'h703: oData <= 1'b1;
            12'h704: oData <= 1'b1;
            12'h705: oData <= 1'b1;
            12'h706: oData <= 1'b1;
            12'h707: oData <= 1'b1;
            12'h708: oData <= 1'b0;
            12'h709: oData <= 1'b0;
            12'h70a: oData <= 1'b0;
            12'h70b: oData <= 1'b0;
            12'h70c: oData <= 1'b0;
            12'h70d: oData <= 1'b0;
            12'h70e: oData <= 1'b0;
            12'h70f: oData <= 1'b0;
            12'h710: oData <= 1'b1;
            12'h711: oData <= 1'b1;
            12'h712: oData <= 1'b1;
            12'h713: oData <= 1'b1;
            12'h714: oData <= 1'b1;
            12'h715: oData <= 1'b1;
            12'h716: oData <= 1'b1;
            12'h717: oData <= 1'b1;
            12'h718: oData <= 1'b0;
            12'h719: oData <= 1'b0;
            12'h71a: oData <= 1'b0;
            12'h71b: oData <= 1'b0;
            12'h71c: oData <= 1'b0;
            12'h71d: oData <= 1'b0;
            12'h71e: oData <= 1'b0;
            12'h71f: oData <= 1'b0;
            12'h720: oData <= 1'b1;
            12'h721: oData <= 1'b1;
            12'h722: oData <= 1'b1;
            12'h723: oData <= 1'b1;
            12'h724: oData <= 1'b1;
            12'h725: oData <= 1'b1;
            12'h726: oData <= 1'b1;
            12'h727: oData <= 1'b0;
            12'h728: oData <= 1'b0;
            12'h729: oData <= 1'b0;
            12'h72a: oData <= 1'b0;
            12'h72b: oData <= 1'b0;
            12'h72c: oData <= 1'b0;
            12'h72d: oData <= 1'b0;
            12'h72e: oData <= 1'b0;
            12'h72f: oData <= 1'b0;
            12'h730: oData <= 1'b1;
            12'h731: oData <= 1'b1;
            12'h732: oData <= 1'b1;
            12'h733: oData <= 1'b1;
            12'h734: oData <= 1'b1;
            12'h735: oData <= 1'b1;
            12'h736: oData <= 1'b1;
            12'h737: oData <= 1'b0;
            12'h738: oData <= 1'b0;
            12'h739: oData <= 1'b0;
            12'h73a: oData <= 1'b0;
            12'h73b: oData <= 1'b0;
            12'h73c: oData <= 1'b0;
            12'h73d: oData <= 1'b0;
            12'h73e: oData <= 1'b0;
            12'h73f: oData <= 1'b0;
            12'h740: oData <= 1'b1;
            12'h741: oData <= 1'b1;
            12'h742: oData <= 1'b1;
            12'h743: oData <= 1'b1;
            12'h744: oData <= 1'b1;
            12'h745: oData <= 1'b1;
            12'h746: oData <= 1'b0;
            12'h747: oData <= 1'b0;
            12'h748: oData <= 1'b0;
            12'h749: oData <= 1'b0;
            12'h74a: oData <= 1'b0;
            12'h74b: oData <= 1'b0;
            12'h74c: oData <= 1'b0;
            12'h74d: oData <= 1'b0;
            12'h74e: oData <= 1'b0;
            12'h74f: oData <= 1'b0;
            12'h750: oData <= 1'b1;
            12'h751: oData <= 1'b1;
            12'h752: oData <= 1'b1;
            12'h753: oData <= 1'b1;
            12'h754: oData <= 1'b1;
            12'h755: oData <= 1'b0;
            12'h756: oData <= 1'b0;
            12'h757: oData <= 1'b0;
            12'h758: oData <= 1'b0;
            12'h759: oData <= 1'b0;
            12'h75a: oData <= 1'b0;
            12'h75b: oData <= 1'b0;
            12'h75c: oData <= 1'b0;
            12'h75d: oData <= 1'b0;
            12'h75e: oData <= 1'b0;
            12'h75f: oData <= 1'b0;
            12'h760: oData <= 1'b1;
            12'h761: oData <= 1'b1;
            12'h762: oData <= 1'b1;
            12'h763: oData <= 1'b1;
            12'h764: oData <= 1'b0;
            12'h765: oData <= 1'b0;
            12'h766: oData <= 1'b0;
            12'h767: oData <= 1'b0;
            12'h768: oData <= 1'b0;
            12'h769: oData <= 1'b0;
            12'h76a: oData <= 1'b0;
            12'h76b: oData <= 1'b0;
            12'h76c: oData <= 1'b0;
            12'h76d: oData <= 1'b0;
            12'h76e: oData <= 1'b0;
            12'h76f: oData <= 1'b0;
            12'h770: oData <= 1'b1;
            12'h771: oData <= 1'b1;
            12'h772: oData <= 1'b0;
            12'h773: oData <= 1'b0;
            12'h774: oData <= 1'b0;
            12'h775: oData <= 1'b0;
            12'h776: oData <= 1'b0;
            12'h777: oData <= 1'b0;
            12'h778: oData <= 1'b0;
            12'h779: oData <= 1'b0;
            12'h77a: oData <= 1'b0;
            12'h77b: oData <= 1'b0;
            12'h77c: oData <= 1'b0;
            12'h77d: oData <= 1'b0;
            12'h77e: oData <= 1'b0;
            12'h77f: oData <= 1'b0;
            12'h780: oData <= 1'b0;
            12'h781: oData <= 1'b0;
            12'h782: oData <= 1'b0;
            12'h783: oData <= 1'b0;
            12'h784: oData <= 1'b0;
            12'h785: oData <= 1'b0;
            12'h786: oData <= 1'b0;
            12'h787: oData <= 1'b0;
            12'h788: oData <= 1'b0;
            12'h789: oData <= 1'b0;
            12'h78a: oData <= 1'b0;
            12'h78b: oData <= 1'b0;
            12'h78c: oData <= 1'b0;
            12'h78d: oData <= 1'b0;
            12'h78e: oData <= 1'b0;
            12'h78f: oData <= 1'b0;
            12'h790: oData <= 1'b0;
            12'h791: oData <= 1'b0;
            12'h792: oData <= 1'b0;
            12'h793: oData <= 1'b0;
            12'h794: oData <= 1'b0;
            12'h795: oData <= 1'b0;
            12'h796: oData <= 1'b0;
            12'h797: oData <= 1'b0;
            12'h798: oData <= 1'b0;
            12'h799: oData <= 1'b0;
            12'h79a: oData <= 1'b0;
            12'h79b: oData <= 1'b0;
            12'h79c: oData <= 1'b0;
            12'h79d: oData <= 1'b0;
            12'h79e: oData <= 1'b0;
            12'h79f: oData <= 1'b0;
            12'h7a0: oData <= 1'b0;
            12'h7a1: oData <= 1'b0;
            12'h7a2: oData <= 1'b0;
            12'h7a3: oData <= 1'b0;
            12'h7a4: oData <= 1'b0;
            12'h7a5: oData <= 1'b0;
            12'h7a6: oData <= 1'b0;
            12'h7a7: oData <= 1'b0;
            12'h7a8: oData <= 1'b0;
            12'h7a9: oData <= 1'b0;
            12'h7aa: oData <= 1'b0;
            12'h7ab: oData <= 1'b0;
            12'h7ac: oData <= 1'b0;
            12'h7ad: oData <= 1'b0;
            12'h7ae: oData <= 1'b0;
            12'h7af: oData <= 1'b0;
            12'h7b0: oData <= 1'b0;
            12'h7b1: oData <= 1'b0;
            12'h7b2: oData <= 1'b0;
            12'h7b3: oData <= 1'b0;
            12'h7b4: oData <= 1'b0;
            12'h7b5: oData <= 1'b0;
            12'h7b6: oData <= 1'b0;
            12'h7b7: oData <= 1'b0;
            12'h7b8: oData <= 1'b0;
            12'h7b9: oData <= 1'b0;
            12'h7ba: oData <= 1'b0;
            12'h7bb: oData <= 1'b0;
            12'h7bc: oData <= 1'b0;
            12'h7bd: oData <= 1'b0;
            12'h7be: oData <= 1'b0;
            12'h7bf: oData <= 1'b0;
            12'h7c0: oData <= 1'b0;
            12'h7c1: oData <= 1'b0;
            12'h7c2: oData <= 1'b0;
            12'h7c3: oData <= 1'b0;
            12'h7c4: oData <= 1'b0;
            12'h7c5: oData <= 1'b0;
            12'h7c6: oData <= 1'b0;
            12'h7c7: oData <= 1'b0;
            12'h7c8: oData <= 1'b0;
            12'h7c9: oData <= 1'b0;
            12'h7ca: oData <= 1'b0;
            12'h7cb: oData <= 1'b0;
            12'h7cc: oData <= 1'b0;
            12'h7cd: oData <= 1'b0;
            12'h7ce: oData <= 1'b0;
            12'h7cf: oData <= 1'b0;
            12'h7d0: oData <= 1'b0;
            12'h7d1: oData <= 1'b0;
            12'h7d2: oData <= 1'b0;
            12'h7d3: oData <= 1'b0;
            12'h7d4: oData <= 1'b0;
            12'h7d5: oData <= 1'b0;
            12'h7d6: oData <= 1'b0;
            12'h7d7: oData <= 1'b0;
            12'h7d8: oData <= 1'b0;
            12'h7d9: oData <= 1'b0;
            12'h7da: oData <= 1'b0;
            12'h7db: oData <= 1'b0;
            12'h7dc: oData <= 1'b0;
            12'h7dd: oData <= 1'b0;
            12'h7de: oData <= 1'b0;
            12'h7df: oData <= 1'b0;
            12'h7e0: oData <= 1'b0;
            12'h7e1: oData <= 1'b0;
            12'h7e2: oData <= 1'b0;
            12'h7e3: oData <= 1'b0;
            12'h7e4: oData <= 1'b0;
            12'h7e5: oData <= 1'b0;
            12'h7e6: oData <= 1'b0;
            12'h7e7: oData <= 1'b0;
            12'h7e8: oData <= 1'b0;
            12'h7e9: oData <= 1'b0;
            12'h7ea: oData <= 1'b0;
            12'h7eb: oData <= 1'b0;
            12'h7ec: oData <= 1'b0;
            12'h7ed: oData <= 1'b0;
            12'h7ee: oData <= 1'b0;
            12'h7ef: oData <= 1'b0;
            12'h7f0: oData <= 1'b0;
            12'h7f1: oData <= 1'b0;
            12'h7f2: oData <= 1'b0;
            12'h7f3: oData <= 1'b0;
            12'h7f4: oData <= 1'b0;
            12'h7f5: oData <= 1'b0;
            12'h7f6: oData <= 1'b0;
            12'h7f7: oData <= 1'b0;
            12'h7f8: oData <= 1'b0;
            12'h7f9: oData <= 1'b0;
            12'h7fa: oData <= 1'b0;
            12'h7fb: oData <= 1'b0;
            12'h7fc: oData <= 1'b0;
            12'h7fd: oData <= 1'b0;
            12'h7fe: oData <= 1'b0;
            12'h7ff: oData <= 1'b0;
            12'h800: oData <= 1'b1;
            12'h801: oData <= 1'b1;
            12'h802: oData <= 1'b1;
            12'h803: oData <= 1'b1;
            12'h804: oData <= 1'b1;
            12'h805: oData <= 1'b1;
            12'h806: oData <= 1'b1;
            12'h807: oData <= 1'b1;
            12'h808: oData <= 1'b1;
            12'h809: oData <= 1'b0;
            12'h80a: oData <= 1'b0;
            12'h80b: oData <= 1'b0;
            12'h80c: oData <= 1'b0;
            12'h80d: oData <= 1'b0;
            12'h80e: oData <= 1'b0;
            12'h80f: oData <= 1'b0;
            12'h810: oData <= 1'b1;
            12'h811: oData <= 1'b1;
            12'h812: oData <= 1'b1;
            12'h813: oData <= 1'b1;
            12'h814: oData <= 1'b1;
            12'h815: oData <= 1'b1;
            12'h816: oData <= 1'b1;
            12'h817: oData <= 1'b1;
            12'h818: oData <= 1'b1;
            12'h819: oData <= 1'b0;
            12'h81a: oData <= 1'b0;
            12'h81b: oData <= 1'b0;
            12'h81c: oData <= 1'b0;
            12'h81d: oData <= 1'b0;
            12'h81e: oData <= 1'b0;
            12'h81f: oData <= 1'b0;
            12'h820: oData <= 1'b1;
            12'h821: oData <= 1'b1;
            12'h822: oData <= 1'b1;
            12'h823: oData <= 1'b1;
            12'h824: oData <= 1'b1;
            12'h825: oData <= 1'b1;
            12'h826: oData <= 1'b1;
            12'h827: oData <= 1'b1;
            12'h828: oData <= 1'b1;
            12'h829: oData <= 1'b0;
            12'h82a: oData <= 1'b0;
            12'h82b: oData <= 1'b0;
            12'h82c: oData <= 1'b0;
            12'h82d: oData <= 1'b0;
            12'h82e: oData <= 1'b0;
            12'h82f: oData <= 1'b0;
            12'h830: oData <= 1'b1;
            12'h831: oData <= 1'b1;
            12'h832: oData <= 1'b1;
            12'h833: oData <= 1'b1;
            12'h834: oData <= 1'b1;
            12'h835: oData <= 1'b1;
            12'h836: oData <= 1'b1;
            12'h837: oData <= 1'b1;
            12'h838: oData <= 1'b0;
            12'h839: oData <= 1'b0;
            12'h83a: oData <= 1'b0;
            12'h83b: oData <= 1'b0;
            12'h83c: oData <= 1'b0;
            12'h83d: oData <= 1'b0;
            12'h83e: oData <= 1'b0;
            12'h83f: oData <= 1'b0;
            12'h840: oData <= 1'b1;
            12'h841: oData <= 1'b1;
            12'h842: oData <= 1'b1;
            12'h843: oData <= 1'b1;
            12'h844: oData <= 1'b1;
            12'h845: oData <= 1'b1;
            12'h846: oData <= 1'b1;
            12'h847: oData <= 1'b1;
            12'h848: oData <= 1'b0;
            12'h849: oData <= 1'b0;
            12'h84a: oData <= 1'b0;
            12'h84b: oData <= 1'b0;
            12'h84c: oData <= 1'b0;
            12'h84d: oData <= 1'b0;
            12'h84e: oData <= 1'b0;
            12'h84f: oData <= 1'b0;
            12'h850: oData <= 1'b1;
            12'h851: oData <= 1'b1;
            12'h852: oData <= 1'b1;
            12'h853: oData <= 1'b1;
            12'h854: oData <= 1'b1;
            12'h855: oData <= 1'b1;
            12'h856: oData <= 1'b1;
            12'h857: oData <= 1'b0;
            12'h858: oData <= 1'b0;
            12'h859: oData <= 1'b0;
            12'h85a: oData <= 1'b0;
            12'h85b: oData <= 1'b0;
            12'h85c: oData <= 1'b0;
            12'h85d: oData <= 1'b0;
            12'h85e: oData <= 1'b0;
            12'h85f: oData <= 1'b0;
            12'h860: oData <= 1'b1;
            12'h861: oData <= 1'b1;
            12'h862: oData <= 1'b1;
            12'h863: oData <= 1'b1;
            12'h864: oData <= 1'b1;
            12'h865: oData <= 1'b1;
            12'h866: oData <= 1'b0;
            12'h867: oData <= 1'b0;
            12'h868: oData <= 1'b0;
            12'h869: oData <= 1'b0;
            12'h86a: oData <= 1'b0;
            12'h86b: oData <= 1'b0;
            12'h86c: oData <= 1'b0;
            12'h86d: oData <= 1'b0;
            12'h86e: oData <= 1'b0;
            12'h86f: oData <= 1'b0;
            12'h870: oData <= 1'b1;
            12'h871: oData <= 1'b1;
            12'h872: oData <= 1'b1;
            12'h873: oData <= 1'b1;
            12'h874: oData <= 1'b1;
            12'h875: oData <= 1'b0;
            12'h876: oData <= 1'b0;
            12'h877: oData <= 1'b0;
            12'h878: oData <= 1'b0;
            12'h879: oData <= 1'b0;
            12'h87a: oData <= 1'b0;
            12'h87b: oData <= 1'b0;
            12'h87c: oData <= 1'b0;
            12'h87d: oData <= 1'b0;
            12'h87e: oData <= 1'b0;
            12'h87f: oData <= 1'b0;
            12'h880: oData <= 1'b1;
            12'h881: oData <= 1'b1;
            12'h882: oData <= 1'b1;
            12'h883: oData <= 1'b0;
            12'h884: oData <= 1'b0;
            12'h885: oData <= 1'b0;
            12'h886: oData <= 1'b0;
            12'h887: oData <= 1'b0;
            12'h888: oData <= 1'b0;
            12'h889: oData <= 1'b0;
            12'h88a: oData <= 1'b0;
            12'h88b: oData <= 1'b0;
            12'h88c: oData <= 1'b0;
            12'h88d: oData <= 1'b0;
            12'h88e: oData <= 1'b0;
            12'h88f: oData <= 1'b0;
            12'h890: oData <= 1'b0;
            12'h891: oData <= 1'b0;
            12'h892: oData <= 1'b0;
            12'h893: oData <= 1'b0;
            12'h894: oData <= 1'b0;
            12'h895: oData <= 1'b0;
            12'h896: oData <= 1'b0;
            12'h897: oData <= 1'b0;
            12'h898: oData <= 1'b0;
            12'h899: oData <= 1'b0;
            12'h89a: oData <= 1'b0;
            12'h89b: oData <= 1'b0;
            12'h89c: oData <= 1'b0;
            12'h89d: oData <= 1'b0;
            12'h89e: oData <= 1'b0;
            12'h89f: oData <= 1'b0;
            12'h8a0: oData <= 1'b0;
            12'h8a1: oData <= 1'b0;
            12'h8a2: oData <= 1'b0;
            12'h8a3: oData <= 1'b0;
            12'h8a4: oData <= 1'b0;
            12'h8a5: oData <= 1'b0;
            12'h8a6: oData <= 1'b0;
            12'h8a7: oData <= 1'b0;
            12'h8a8: oData <= 1'b0;
            12'h8a9: oData <= 1'b0;
            12'h8aa: oData <= 1'b0;
            12'h8ab: oData <= 1'b0;
            12'h8ac: oData <= 1'b0;
            12'h8ad: oData <= 1'b0;
            12'h8ae: oData <= 1'b0;
            12'h8af: oData <= 1'b0;
            12'h8b0: oData <= 1'b0;
            12'h8b1: oData <= 1'b0;
            12'h8b2: oData <= 1'b0;
            12'h8b3: oData <= 1'b0;
            12'h8b4: oData <= 1'b0;
            12'h8b5: oData <= 1'b0;
            12'h8b6: oData <= 1'b0;
            12'h8b7: oData <= 1'b0;
            12'h8b8: oData <= 1'b0;
            12'h8b9: oData <= 1'b0;
            12'h8ba: oData <= 1'b0;
            12'h8bb: oData <= 1'b0;
            12'h8bc: oData <= 1'b0;
            12'h8bd: oData <= 1'b0;
            12'h8be: oData <= 1'b0;
            12'h8bf: oData <= 1'b0;
            12'h8c0: oData <= 1'b0;
            12'h8c1: oData <= 1'b0;
            12'h8c2: oData <= 1'b0;
            12'h8c3: oData <= 1'b0;
            12'h8c4: oData <= 1'b0;
            12'h8c5: oData <= 1'b0;
            12'h8c6: oData <= 1'b0;
            12'h8c7: oData <= 1'b0;
            12'h8c8: oData <= 1'b0;
            12'h8c9: oData <= 1'b0;
            12'h8ca: oData <= 1'b0;
            12'h8cb: oData <= 1'b0;
            12'h8cc: oData <= 1'b0;
            12'h8cd: oData <= 1'b0;
            12'h8ce: oData <= 1'b0;
            12'h8cf: oData <= 1'b0;
            12'h8d0: oData <= 1'b0;
            12'h8d1: oData <= 1'b0;
            12'h8d2: oData <= 1'b0;
            12'h8d3: oData <= 1'b0;
            12'h8d4: oData <= 1'b0;
            12'h8d5: oData <= 1'b0;
            12'h8d6: oData <= 1'b0;
            12'h8d7: oData <= 1'b0;
            12'h8d8: oData <= 1'b0;
            12'h8d9: oData <= 1'b0;
            12'h8da: oData <= 1'b0;
            12'h8db: oData <= 1'b0;
            12'h8dc: oData <= 1'b0;
            12'h8dd: oData <= 1'b0;
            12'h8de: oData <= 1'b0;
            12'h8df: oData <= 1'b0;
            12'h8e0: oData <= 1'b0;
            12'h8e1: oData <= 1'b0;
            12'h8e2: oData <= 1'b0;
            12'h8e3: oData <= 1'b0;
            12'h8e4: oData <= 1'b0;
            12'h8e5: oData <= 1'b0;
            12'h8e6: oData <= 1'b0;
            12'h8e7: oData <= 1'b0;
            12'h8e8: oData <= 1'b0;
            12'h8e9: oData <= 1'b0;
            12'h8ea: oData <= 1'b0;
            12'h8eb: oData <= 1'b0;
            12'h8ec: oData <= 1'b0;
            12'h8ed: oData <= 1'b0;
            12'h8ee: oData <= 1'b0;
            12'h8ef: oData <= 1'b0;
            12'h8f0: oData <= 1'b0;
            12'h8f1: oData <= 1'b0;
            12'h8f2: oData <= 1'b0;
            12'h8f3: oData <= 1'b0;
            12'h8f4: oData <= 1'b0;
            12'h8f5: oData <= 1'b0;
            12'h8f6: oData <= 1'b0;
            12'h8f7: oData <= 1'b0;
            12'h8f8: oData <= 1'b0;
            12'h8f9: oData <= 1'b0;
            12'h8fa: oData <= 1'b0;
            12'h8fb: oData <= 1'b0;
            12'h8fc: oData <= 1'b0;
            12'h8fd: oData <= 1'b0;
            12'h8fe: oData <= 1'b0;
            12'h8ff: oData <= 1'b0;
            12'h900: oData <= 1'b1;
            12'h901: oData <= 1'b1;
            12'h902: oData <= 1'b1;
            12'h903: oData <= 1'b1;
            12'h904: oData <= 1'b1;
            12'h905: oData <= 1'b1;
            12'h906: oData <= 1'b1;
            12'h907: oData <= 1'b1;
            12'h908: oData <= 1'b1;
            12'h909: oData <= 1'b1;
            12'h90a: oData <= 1'b0;
            12'h90b: oData <= 1'b0;
            12'h90c: oData <= 1'b0;
            12'h90d: oData <= 1'b0;
            12'h90e: oData <= 1'b0;
            12'h90f: oData <= 1'b0;
            12'h910: oData <= 1'b1;
            12'h911: oData <= 1'b1;
            12'h912: oData <= 1'b1;
            12'h913: oData <= 1'b1;
            12'h914: oData <= 1'b1;
            12'h915: oData <= 1'b1;
            12'h916: oData <= 1'b1;
            12'h917: oData <= 1'b1;
            12'h918: oData <= 1'b1;
            12'h919: oData <= 1'b1;
            12'h91a: oData <= 1'b0;
            12'h91b: oData <= 1'b0;
            12'h91c: oData <= 1'b0;
            12'h91d: oData <= 1'b0;
            12'h91e: oData <= 1'b0;
            12'h91f: oData <= 1'b0;
            12'h920: oData <= 1'b1;
            12'h921: oData <= 1'b1;
            12'h922: oData <= 1'b1;
            12'h923: oData <= 1'b1;
            12'h924: oData <= 1'b1;
            12'h925: oData <= 1'b1;
            12'h926: oData <= 1'b1;
            12'h927: oData <= 1'b1;
            12'h928: oData <= 1'b1;
            12'h929: oData <= 1'b1;
            12'h92a: oData <= 1'b0;
            12'h92b: oData <= 1'b0;
            12'h92c: oData <= 1'b0;
            12'h92d: oData <= 1'b0;
            12'h92e: oData <= 1'b0;
            12'h92f: oData <= 1'b0;
            12'h930: oData <= 1'b1;
            12'h931: oData <= 1'b1;
            12'h932: oData <= 1'b1;
            12'h933: oData <= 1'b1;
            12'h934: oData <= 1'b1;
            12'h935: oData <= 1'b1;
            12'h936: oData <= 1'b1;
            12'h937: oData <= 1'b1;
            12'h938: oData <= 1'b1;
            12'h939: oData <= 1'b0;
            12'h93a: oData <= 1'b0;
            12'h93b: oData <= 1'b0;
            12'h93c: oData <= 1'b0;
            12'h93d: oData <= 1'b0;
            12'h93e: oData <= 1'b0;
            12'h93f: oData <= 1'b0;
            12'h940: oData <= 1'b1;
            12'h941: oData <= 1'b1;
            12'h942: oData <= 1'b1;
            12'h943: oData <= 1'b1;
            12'h944: oData <= 1'b1;
            12'h945: oData <= 1'b1;
            12'h946: oData <= 1'b1;
            12'h947: oData <= 1'b1;
            12'h948: oData <= 1'b1;
            12'h949: oData <= 1'b0;
            12'h94a: oData <= 1'b0;
            12'h94b: oData <= 1'b0;
            12'h94c: oData <= 1'b0;
            12'h94d: oData <= 1'b0;
            12'h94e: oData <= 1'b0;
            12'h94f: oData <= 1'b0;
            12'h950: oData <= 1'b1;
            12'h951: oData <= 1'b1;
            12'h952: oData <= 1'b1;
            12'h953: oData <= 1'b1;
            12'h954: oData <= 1'b1;
            12'h955: oData <= 1'b1;
            12'h956: oData <= 1'b1;
            12'h957: oData <= 1'b1;
            12'h958: oData <= 1'b1;
            12'h959: oData <= 1'b0;
            12'h95a: oData <= 1'b0;
            12'h95b: oData <= 1'b0;
            12'h95c: oData <= 1'b0;
            12'h95d: oData <= 1'b0;
            12'h95e: oData <= 1'b0;
            12'h95f: oData <= 1'b0;
            12'h960: oData <= 1'b1;
            12'h961: oData <= 1'b1;
            12'h962: oData <= 1'b1;
            12'h963: oData <= 1'b1;
            12'h964: oData <= 1'b1;
            12'h965: oData <= 1'b1;
            12'h966: oData <= 1'b1;
            12'h967: oData <= 1'b1;
            12'h968: oData <= 1'b0;
            12'h969: oData <= 1'b0;
            12'h96a: oData <= 1'b0;
            12'h96b: oData <= 1'b0;
            12'h96c: oData <= 1'b0;
            12'h96d: oData <= 1'b0;
            12'h96e: oData <= 1'b0;
            12'h96f: oData <= 1'b0;
            12'h970: oData <= 1'b1;
            12'h971: oData <= 1'b1;
            12'h972: oData <= 1'b1;
            12'h973: oData <= 1'b1;
            12'h974: oData <= 1'b1;
            12'h975: oData <= 1'b1;
            12'h976: oData <= 1'b1;
            12'h977: oData <= 1'b0;
            12'h978: oData <= 1'b0;
            12'h979: oData <= 1'b0;
            12'h97a: oData <= 1'b0;
            12'h97b: oData <= 1'b0;
            12'h97c: oData <= 1'b0;
            12'h97d: oData <= 1'b0;
            12'h97e: oData <= 1'b0;
            12'h97f: oData <= 1'b0;
            12'h980: oData <= 1'b1;
            12'h981: oData <= 1'b1;
            12'h982: oData <= 1'b1;
            12'h983: oData <= 1'b1;
            12'h984: oData <= 1'b1;
            12'h985: oData <= 1'b1;
            12'h986: oData <= 1'b0;
            12'h987: oData <= 1'b0;
            12'h988: oData <= 1'b0;
            12'h989: oData <= 1'b0;
            12'h98a: oData <= 1'b0;
            12'h98b: oData <= 1'b0;
            12'h98c: oData <= 1'b0;
            12'h98d: oData <= 1'b0;
            12'h98e: oData <= 1'b0;
            12'h98f: oData <= 1'b0;
            12'h990: oData <= 1'b1;
            12'h991: oData <= 1'b1;
            12'h992: oData <= 1'b1;
            12'h993: oData <= 1'b0;
            12'h994: oData <= 1'b0;
            12'h995: oData <= 1'b0;
            12'h996: oData <= 1'b0;
            12'h997: oData <= 1'b0;
            12'h998: oData <= 1'b0;
            12'h999: oData <= 1'b0;
            12'h99a: oData <= 1'b0;
            12'h99b: oData <= 1'b0;
            12'h99c: oData <= 1'b0;
            12'h99d: oData <= 1'b0;
            12'h99e: oData <= 1'b0;
            12'h99f: oData <= 1'b0;
            12'h9a0: oData <= 1'b0;
            12'h9a1: oData <= 1'b0;
            12'h9a2: oData <= 1'b0;
            12'h9a3: oData <= 1'b0;
            12'h9a4: oData <= 1'b0;
            12'h9a5: oData <= 1'b0;
            12'h9a6: oData <= 1'b0;
            12'h9a7: oData <= 1'b0;
            12'h9a8: oData <= 1'b0;
            12'h9a9: oData <= 1'b0;
            12'h9aa: oData <= 1'b0;
            12'h9ab: oData <= 1'b0;
            12'h9ac: oData <= 1'b0;
            12'h9ad: oData <= 1'b0;
            12'h9ae: oData <= 1'b0;
            12'h9af: oData <= 1'b0;
            12'h9b0: oData <= 1'b0;
            12'h9b1: oData <= 1'b0;
            12'h9b2: oData <= 1'b0;
            12'h9b3: oData <= 1'b0;
            12'h9b4: oData <= 1'b0;
            12'h9b5: oData <= 1'b0;
            12'h9b6: oData <= 1'b0;
            12'h9b7: oData <= 1'b0;
            12'h9b8: oData <= 1'b0;
            12'h9b9: oData <= 1'b0;
            12'h9ba: oData <= 1'b0;
            12'h9bb: oData <= 1'b0;
            12'h9bc: oData <= 1'b0;
            12'h9bd: oData <= 1'b0;
            12'h9be: oData <= 1'b0;
            12'h9bf: oData <= 1'b0;
            12'h9c0: oData <= 1'b0;
            12'h9c1: oData <= 1'b0;
            12'h9c2: oData <= 1'b0;
            12'h9c3: oData <= 1'b0;
            12'h9c4: oData <= 1'b0;
            12'h9c5: oData <= 1'b0;
            12'h9c6: oData <= 1'b0;
            12'h9c7: oData <= 1'b0;
            12'h9c8: oData <= 1'b0;
            12'h9c9: oData <= 1'b0;
            12'h9ca: oData <= 1'b0;
            12'h9cb: oData <= 1'b0;
            12'h9cc: oData <= 1'b0;
            12'h9cd: oData <= 1'b0;
            12'h9ce: oData <= 1'b0;
            12'h9cf: oData <= 1'b0;
            12'h9d0: oData <= 1'b0;
            12'h9d1: oData <= 1'b0;
            12'h9d2: oData <= 1'b0;
            12'h9d3: oData <= 1'b0;
            12'h9d4: oData <= 1'b0;
            12'h9d5: oData <= 1'b0;
            12'h9d6: oData <= 1'b0;
            12'h9d7: oData <= 1'b0;
            12'h9d8: oData <= 1'b0;
            12'h9d9: oData <= 1'b0;
            12'h9da: oData <= 1'b0;
            12'h9db: oData <= 1'b0;
            12'h9dc: oData <= 1'b0;
            12'h9dd: oData <= 1'b0;
            12'h9de: oData <= 1'b0;
            12'h9df: oData <= 1'b0;
            12'h9e0: oData <= 1'b0;
            12'h9e1: oData <= 1'b0;
            12'h9e2: oData <= 1'b0;
            12'h9e3: oData <= 1'b0;
            12'h9e4: oData <= 1'b0;
            12'h9e5: oData <= 1'b0;
            12'h9e6: oData <= 1'b0;
            12'h9e7: oData <= 1'b0;
            12'h9e8: oData <= 1'b0;
            12'h9e9: oData <= 1'b0;
            12'h9ea: oData <= 1'b0;
            12'h9eb: oData <= 1'b0;
            12'h9ec: oData <= 1'b0;
            12'h9ed: oData <= 1'b0;
            12'h9ee: oData <= 1'b0;
            12'h9ef: oData <= 1'b0;
            12'h9f0: oData <= 1'b0;
            12'h9f1: oData <= 1'b0;
            12'h9f2: oData <= 1'b0;
            12'h9f3: oData <= 1'b0;
            12'h9f4: oData <= 1'b0;
            12'h9f5: oData <= 1'b0;
            12'h9f6: oData <= 1'b0;
            12'h9f7: oData <= 1'b0;
            12'h9f8: oData <= 1'b0;
            12'h9f9: oData <= 1'b0;
            12'h9fa: oData <= 1'b0;
            12'h9fb: oData <= 1'b0;
            12'h9fc: oData <= 1'b0;
            12'h9fd: oData <= 1'b0;
            12'h9fe: oData <= 1'b0;
            12'h9ff: oData <= 1'b0;
            12'ha00: oData <= 1'b1;
            12'ha01: oData <= 1'b1;
            12'ha02: oData <= 1'b1;
            12'ha03: oData <= 1'b1;
            12'ha04: oData <= 1'b1;
            12'ha05: oData <= 1'b1;
            12'ha06: oData <= 1'b1;
            12'ha07: oData <= 1'b1;
            12'ha08: oData <= 1'b1;
            12'ha09: oData <= 1'b1;
            12'ha0a: oData <= 1'b1;
            12'ha0b: oData <= 1'b0;
            12'ha0c: oData <= 1'b0;
            12'ha0d: oData <= 1'b0;
            12'ha0e: oData <= 1'b0;
            12'ha0f: oData <= 1'b0;
            12'ha10: oData <= 1'b1;
            12'ha11: oData <= 1'b1;
            12'ha12: oData <= 1'b1;
            12'ha13: oData <= 1'b1;
            12'ha14: oData <= 1'b1;
            12'ha15: oData <= 1'b1;
            12'ha16: oData <= 1'b1;
            12'ha17: oData <= 1'b1;
            12'ha18: oData <= 1'b1;
            12'ha19: oData <= 1'b1;
            12'ha1a: oData <= 1'b1;
            12'ha1b: oData <= 1'b0;
            12'ha1c: oData <= 1'b0;
            12'ha1d: oData <= 1'b0;
            12'ha1e: oData <= 1'b0;
            12'ha1f: oData <= 1'b0;
            12'ha20: oData <= 1'b1;
            12'ha21: oData <= 1'b1;
            12'ha22: oData <= 1'b1;
            12'ha23: oData <= 1'b1;
            12'ha24: oData <= 1'b1;
            12'ha25: oData <= 1'b1;
            12'ha26: oData <= 1'b1;
            12'ha27: oData <= 1'b1;
            12'ha28: oData <= 1'b1;
            12'ha29: oData <= 1'b1;
            12'ha2a: oData <= 1'b1;
            12'ha2b: oData <= 1'b0;
            12'ha2c: oData <= 1'b0;
            12'ha2d: oData <= 1'b0;
            12'ha2e: oData <= 1'b0;
            12'ha2f: oData <= 1'b0;
            12'ha30: oData <= 1'b1;
            12'ha31: oData <= 1'b1;
            12'ha32: oData <= 1'b1;
            12'ha33: oData <= 1'b1;
            12'ha34: oData <= 1'b1;
            12'ha35: oData <= 1'b1;
            12'ha36: oData <= 1'b1;
            12'ha37: oData <= 1'b1;
            12'ha38: oData <= 1'b1;
            12'ha39: oData <= 1'b1;
            12'ha3a: oData <= 1'b0;
            12'ha3b: oData <= 1'b0;
            12'ha3c: oData <= 1'b0;
            12'ha3d: oData <= 1'b0;
            12'ha3e: oData <= 1'b0;
            12'ha3f: oData <= 1'b0;
            12'ha40: oData <= 1'b1;
            12'ha41: oData <= 1'b1;
            12'ha42: oData <= 1'b1;
            12'ha43: oData <= 1'b1;
            12'ha44: oData <= 1'b1;
            12'ha45: oData <= 1'b1;
            12'ha46: oData <= 1'b1;
            12'ha47: oData <= 1'b1;
            12'ha48: oData <= 1'b1;
            12'ha49: oData <= 1'b1;
            12'ha4a: oData <= 1'b0;
            12'ha4b: oData <= 1'b0;
            12'ha4c: oData <= 1'b0;
            12'ha4d: oData <= 1'b0;
            12'ha4e: oData <= 1'b0;
            12'ha4f: oData <= 1'b0;
            12'ha50: oData <= 1'b1;
            12'ha51: oData <= 1'b1;
            12'ha52: oData <= 1'b1;
            12'ha53: oData <= 1'b1;
            12'ha54: oData <= 1'b1;
            12'ha55: oData <= 1'b1;
            12'ha56: oData <= 1'b1;
            12'ha57: oData <= 1'b1;
            12'ha58: oData <= 1'b1;
            12'ha59: oData <= 1'b1;
            12'ha5a: oData <= 1'b0;
            12'ha5b: oData <= 1'b0;
            12'ha5c: oData <= 1'b0;
            12'ha5d: oData <= 1'b0;
            12'ha5e: oData <= 1'b0;
            12'ha5f: oData <= 1'b0;
            12'ha60: oData <= 1'b1;
            12'ha61: oData <= 1'b1;
            12'ha62: oData <= 1'b1;
            12'ha63: oData <= 1'b1;
            12'ha64: oData <= 1'b1;
            12'ha65: oData <= 1'b1;
            12'ha66: oData <= 1'b1;
            12'ha67: oData <= 1'b1;
            12'ha68: oData <= 1'b1;
            12'ha69: oData <= 1'b0;
            12'ha6a: oData <= 1'b0;
            12'ha6b: oData <= 1'b0;
            12'ha6c: oData <= 1'b0;
            12'ha6d: oData <= 1'b0;
            12'ha6e: oData <= 1'b0;
            12'ha6f: oData <= 1'b0;
            12'ha70: oData <= 1'b1;
            12'ha71: oData <= 1'b1;
            12'ha72: oData <= 1'b1;
            12'ha73: oData <= 1'b1;
            12'ha74: oData <= 1'b1;
            12'ha75: oData <= 1'b1;
            12'ha76: oData <= 1'b1;
            12'ha77: oData <= 1'b1;
            12'ha78: oData <= 1'b0;
            12'ha79: oData <= 1'b0;
            12'ha7a: oData <= 1'b0;
            12'ha7b: oData <= 1'b0;
            12'ha7c: oData <= 1'b0;
            12'ha7d: oData <= 1'b0;
            12'ha7e: oData <= 1'b0;
            12'ha7f: oData <= 1'b0;
            12'ha80: oData <= 1'b1;
            12'ha81: oData <= 1'b1;
            12'ha82: oData <= 1'b1;
            12'ha83: oData <= 1'b1;
            12'ha84: oData <= 1'b1;
            12'ha85: oData <= 1'b1;
            12'ha86: oData <= 1'b1;
            12'ha87: oData <= 1'b0;
            12'ha88: oData <= 1'b0;
            12'ha89: oData <= 1'b0;
            12'ha8a: oData <= 1'b0;
            12'ha8b: oData <= 1'b0;
            12'ha8c: oData <= 1'b0;
            12'ha8d: oData <= 1'b0;
            12'ha8e: oData <= 1'b0;
            12'ha8f: oData <= 1'b0;
            12'ha90: oData <= 1'b1;
            12'ha91: oData <= 1'b1;
            12'ha92: oData <= 1'b1;
            12'ha93: oData <= 1'b1;
            12'ha94: oData <= 1'b1;
            12'ha95: oData <= 1'b1;
            12'ha96: oData <= 1'b0;
            12'ha97: oData <= 1'b0;
            12'ha98: oData <= 1'b0;
            12'ha99: oData <= 1'b0;
            12'ha9a: oData <= 1'b0;
            12'ha9b: oData <= 1'b0;
            12'ha9c: oData <= 1'b0;
            12'ha9d: oData <= 1'b0;
            12'ha9e: oData <= 1'b0;
            12'ha9f: oData <= 1'b0;
            12'haa0: oData <= 1'b1;
            12'haa1: oData <= 1'b1;
            12'haa2: oData <= 1'b1;
            12'haa3: oData <= 1'b0;
            12'haa4: oData <= 1'b0;
            12'haa5: oData <= 1'b0;
            12'haa6: oData <= 1'b0;
            12'haa7: oData <= 1'b0;
            12'haa8: oData <= 1'b0;
            12'haa9: oData <= 1'b0;
            12'haaa: oData <= 1'b0;
            12'haab: oData <= 1'b0;
            12'haac: oData <= 1'b0;
            12'haad: oData <= 1'b0;
            12'haae: oData <= 1'b0;
            12'haaf: oData <= 1'b0;
            12'hab0: oData <= 1'b0;
            12'hab1: oData <= 1'b0;
            12'hab2: oData <= 1'b0;
            12'hab3: oData <= 1'b0;
            12'hab4: oData <= 1'b0;
            12'hab5: oData <= 1'b0;
            12'hab6: oData <= 1'b0;
            12'hab7: oData <= 1'b0;
            12'hab8: oData <= 1'b0;
            12'hab9: oData <= 1'b0;
            12'haba: oData <= 1'b0;
            12'habb: oData <= 1'b0;
            12'habc: oData <= 1'b0;
            12'habd: oData <= 1'b0;
            12'habe: oData <= 1'b0;
            12'habf: oData <= 1'b0;
            12'hac0: oData <= 1'b0;
            12'hac1: oData <= 1'b0;
            12'hac2: oData <= 1'b0;
            12'hac3: oData <= 1'b0;
            12'hac4: oData <= 1'b0;
            12'hac5: oData <= 1'b0;
            12'hac6: oData <= 1'b0;
            12'hac7: oData <= 1'b0;
            12'hac8: oData <= 1'b0;
            12'hac9: oData <= 1'b0;
            12'haca: oData <= 1'b0;
            12'hacb: oData <= 1'b0;
            12'hacc: oData <= 1'b0;
            12'hacd: oData <= 1'b0;
            12'hace: oData <= 1'b0;
            12'hacf: oData <= 1'b0;
            12'had0: oData <= 1'b0;
            12'had1: oData <= 1'b0;
            12'had2: oData <= 1'b0;
            12'had3: oData <= 1'b0;
            12'had4: oData <= 1'b0;
            12'had5: oData <= 1'b0;
            12'had6: oData <= 1'b0;
            12'had7: oData <= 1'b0;
            12'had8: oData <= 1'b0;
            12'had9: oData <= 1'b0;
            12'hada: oData <= 1'b0;
            12'hadb: oData <= 1'b0;
            12'hadc: oData <= 1'b0;
            12'hadd: oData <= 1'b0;
            12'hade: oData <= 1'b0;
            12'hadf: oData <= 1'b0;
            12'hae0: oData <= 1'b0;
            12'hae1: oData <= 1'b0;
            12'hae2: oData <= 1'b0;
            12'hae3: oData <= 1'b0;
            12'hae4: oData <= 1'b0;
            12'hae5: oData <= 1'b0;
            12'hae6: oData <= 1'b0;
            12'hae7: oData <= 1'b0;
            12'hae8: oData <= 1'b0;
            12'hae9: oData <= 1'b0;
            12'haea: oData <= 1'b0;
            12'haeb: oData <= 1'b0;
            12'haec: oData <= 1'b0;
            12'haed: oData <= 1'b0;
            12'haee: oData <= 1'b0;
            12'haef: oData <= 1'b0;
            12'haf0: oData <= 1'b0;
            12'haf1: oData <= 1'b0;
            12'haf2: oData <= 1'b0;
            12'haf3: oData <= 1'b0;
            12'haf4: oData <= 1'b0;
            12'haf5: oData <= 1'b0;
            12'haf6: oData <= 1'b0;
            12'haf7: oData <= 1'b0;
            12'haf8: oData <= 1'b0;
            12'haf9: oData <= 1'b0;
            12'hafa: oData <= 1'b0;
            12'hafb: oData <= 1'b0;
            12'hafc: oData <= 1'b0;
            12'hafd: oData <= 1'b0;
            12'hafe: oData <= 1'b0;
            12'haff: oData <= 1'b0;
            12'hb00: oData <= 1'b1;
            12'hb01: oData <= 1'b1;
            12'hb02: oData <= 1'b1;
            12'hb03: oData <= 1'b1;
            12'hb04: oData <= 1'b1;
            12'hb05: oData <= 1'b1;
            12'hb06: oData <= 1'b1;
            12'hb07: oData <= 1'b1;
            12'hb08: oData <= 1'b1;
            12'hb09: oData <= 1'b1;
            12'hb0a: oData <= 1'b1;
            12'hb0b: oData <= 1'b1;
            12'hb0c: oData <= 1'b0;
            12'hb0d: oData <= 1'b0;
            12'hb0e: oData <= 1'b0;
            12'hb0f: oData <= 1'b0;
            12'hb10: oData <= 1'b1;
            12'hb11: oData <= 1'b1;
            12'hb12: oData <= 1'b1;
            12'hb13: oData <= 1'b1;
            12'hb14: oData <= 1'b1;
            12'hb15: oData <= 1'b1;
            12'hb16: oData <= 1'b1;
            12'hb17: oData <= 1'b1;
            12'hb18: oData <= 1'b1;
            12'hb19: oData <= 1'b1;
            12'hb1a: oData <= 1'b1;
            12'hb1b: oData <= 1'b1;
            12'hb1c: oData <= 1'b0;
            12'hb1d: oData <= 1'b0;
            12'hb1e: oData <= 1'b0;
            12'hb1f: oData <= 1'b0;
            12'hb20: oData <= 1'b1;
            12'hb21: oData <= 1'b1;
            12'hb22: oData <= 1'b1;
            12'hb23: oData <= 1'b1;
            12'hb24: oData <= 1'b1;
            12'hb25: oData <= 1'b1;
            12'hb26: oData <= 1'b1;
            12'hb27: oData <= 1'b1;
            12'hb28: oData <= 1'b1;
            12'hb29: oData <= 1'b1;
            12'hb2a: oData <= 1'b1;
            12'hb2b: oData <= 1'b1;
            12'hb2c: oData <= 1'b0;
            12'hb2d: oData <= 1'b0;
            12'hb2e: oData <= 1'b0;
            12'hb2f: oData <= 1'b0;
            12'hb30: oData <= 1'b1;
            12'hb31: oData <= 1'b1;
            12'hb32: oData <= 1'b1;
            12'hb33: oData <= 1'b1;
            12'hb34: oData <= 1'b1;
            12'hb35: oData <= 1'b1;
            12'hb36: oData <= 1'b1;
            12'hb37: oData <= 1'b1;
            12'hb38: oData <= 1'b1;
            12'hb39: oData <= 1'b1;
            12'hb3a: oData <= 1'b1;
            12'hb3b: oData <= 1'b0;
            12'hb3c: oData <= 1'b0;
            12'hb3d: oData <= 1'b0;
            12'hb3e: oData <= 1'b0;
            12'hb3f: oData <= 1'b0;
            12'hb40: oData <= 1'b1;
            12'hb41: oData <= 1'b1;
            12'hb42: oData <= 1'b1;
            12'hb43: oData <= 1'b1;
            12'hb44: oData <= 1'b1;
            12'hb45: oData <= 1'b1;
            12'hb46: oData <= 1'b1;
            12'hb47: oData <= 1'b1;
            12'hb48: oData <= 1'b1;
            12'hb49: oData <= 1'b1;
            12'hb4a: oData <= 1'b1;
            12'hb4b: oData <= 1'b0;
            12'hb4c: oData <= 1'b0;
            12'hb4d: oData <= 1'b0;
            12'hb4e: oData <= 1'b0;
            12'hb4f: oData <= 1'b0;
            12'hb50: oData <= 1'b1;
            12'hb51: oData <= 1'b1;
            12'hb52: oData <= 1'b1;
            12'hb53: oData <= 1'b1;
            12'hb54: oData <= 1'b1;
            12'hb55: oData <= 1'b1;
            12'hb56: oData <= 1'b1;
            12'hb57: oData <= 1'b1;
            12'hb58: oData <= 1'b1;
            12'hb59: oData <= 1'b1;
            12'hb5a: oData <= 1'b1;
            12'hb5b: oData <= 1'b0;
            12'hb5c: oData <= 1'b0;
            12'hb5d: oData <= 1'b0;
            12'hb5e: oData <= 1'b0;
            12'hb5f: oData <= 1'b0;
            12'hb60: oData <= 1'b1;
            12'hb61: oData <= 1'b1;
            12'hb62: oData <= 1'b1;
            12'hb63: oData <= 1'b1;
            12'hb64: oData <= 1'b1;
            12'hb65: oData <= 1'b1;
            12'hb66: oData <= 1'b1;
            12'hb67: oData <= 1'b1;
            12'hb68: oData <= 1'b1;
            12'hb69: oData <= 1'b1;
            12'hb6a: oData <= 1'b0;
            12'hb6b: oData <= 1'b0;
            12'hb6c: oData <= 1'b0;
            12'hb6d: oData <= 1'b0;
            12'hb6e: oData <= 1'b0;
            12'hb6f: oData <= 1'b0;
            12'hb70: oData <= 1'b1;
            12'hb71: oData <= 1'b1;
            12'hb72: oData <= 1'b1;
            12'hb73: oData <= 1'b1;
            12'hb74: oData <= 1'b1;
            12'hb75: oData <= 1'b1;
            12'hb76: oData <= 1'b1;
            12'hb77: oData <= 1'b1;
            12'hb78: oData <= 1'b1;
            12'hb79: oData <= 1'b1;
            12'hb7a: oData <= 1'b0;
            12'hb7b: oData <= 1'b0;
            12'hb7c: oData <= 1'b0;
            12'hb7d: oData <= 1'b0;
            12'hb7e: oData <= 1'b0;
            12'hb7f: oData <= 1'b0;
            12'hb80: oData <= 1'b1;
            12'hb81: oData <= 1'b1;
            12'hb82: oData <= 1'b1;
            12'hb83: oData <= 1'b1;
            12'hb84: oData <= 1'b1;
            12'hb85: oData <= 1'b1;
            12'hb86: oData <= 1'b1;
            12'hb87: oData <= 1'b1;
            12'hb88: oData <= 1'b1;
            12'hb89: oData <= 1'b0;
            12'hb8a: oData <= 1'b0;
            12'hb8b: oData <= 1'b0;
            12'hb8c: oData <= 1'b0;
            12'hb8d: oData <= 1'b0;
            12'hb8e: oData <= 1'b0;
            12'hb8f: oData <= 1'b0;
            12'hb90: oData <= 1'b1;
            12'hb91: oData <= 1'b1;
            12'hb92: oData <= 1'b1;
            12'hb93: oData <= 1'b1;
            12'hb94: oData <= 1'b1;
            12'hb95: oData <= 1'b1;
            12'hb96: oData <= 1'b1;
            12'hb97: oData <= 1'b1;
            12'hb98: oData <= 1'b0;
            12'hb99: oData <= 1'b0;
            12'hb9a: oData <= 1'b0;
            12'hb9b: oData <= 1'b0;
            12'hb9c: oData <= 1'b0;
            12'hb9d: oData <= 1'b0;
            12'hb9e: oData <= 1'b0;
            12'hb9f: oData <= 1'b0;
            12'hba0: oData <= 1'b1;
            12'hba1: oData <= 1'b1;
            12'hba2: oData <= 1'b1;
            12'hba3: oData <= 1'b1;
            12'hba4: oData <= 1'b1;
            12'hba5: oData <= 1'b1;
            12'hba6: oData <= 1'b0;
            12'hba7: oData <= 1'b0;
            12'hba8: oData <= 1'b0;
            12'hba9: oData <= 1'b0;
            12'hbaa: oData <= 1'b0;
            12'hbab: oData <= 1'b0;
            12'hbac: oData <= 1'b0;
            12'hbad: oData <= 1'b0;
            12'hbae: oData <= 1'b0;
            12'hbaf: oData <= 1'b0;
            12'hbb0: oData <= 1'b1;
            12'hbb1: oData <= 1'b1;
            12'hbb2: oData <= 1'b1;
            12'hbb3: oData <= 1'b0;
            12'hbb4: oData <= 1'b0;
            12'hbb5: oData <= 1'b0;
            12'hbb6: oData <= 1'b0;
            12'hbb7: oData <= 1'b0;
            12'hbb8: oData <= 1'b0;
            12'hbb9: oData <= 1'b0;
            12'hbba: oData <= 1'b0;
            12'hbbb: oData <= 1'b0;
            12'hbbc: oData <= 1'b0;
            12'hbbd: oData <= 1'b0;
            12'hbbe: oData <= 1'b0;
            12'hbbf: oData <= 1'b0;
            12'hbc0: oData <= 1'b0;
            12'hbc1: oData <= 1'b0;
            12'hbc2: oData <= 1'b0;
            12'hbc3: oData <= 1'b0;
            12'hbc4: oData <= 1'b0;
            12'hbc5: oData <= 1'b0;
            12'hbc6: oData <= 1'b0;
            12'hbc7: oData <= 1'b0;
            12'hbc8: oData <= 1'b0;
            12'hbc9: oData <= 1'b0;
            12'hbca: oData <= 1'b0;
            12'hbcb: oData <= 1'b0;
            12'hbcc: oData <= 1'b0;
            12'hbcd: oData <= 1'b0;
            12'hbce: oData <= 1'b0;
            12'hbcf: oData <= 1'b0;
            12'hbd0: oData <= 1'b0;
            12'hbd1: oData <= 1'b0;
            12'hbd2: oData <= 1'b0;
            12'hbd3: oData <= 1'b0;
            12'hbd4: oData <= 1'b0;
            12'hbd5: oData <= 1'b0;
            12'hbd6: oData <= 1'b0;
            12'hbd7: oData <= 1'b0;
            12'hbd8: oData <= 1'b0;
            12'hbd9: oData <= 1'b0;
            12'hbda: oData <= 1'b0;
            12'hbdb: oData <= 1'b0;
            12'hbdc: oData <= 1'b0;
            12'hbdd: oData <= 1'b0;
            12'hbde: oData <= 1'b0;
            12'hbdf: oData <= 1'b0;
            12'hbe0: oData <= 1'b0;
            12'hbe1: oData <= 1'b0;
            12'hbe2: oData <= 1'b0;
            12'hbe3: oData <= 1'b0;
            12'hbe4: oData <= 1'b0;
            12'hbe5: oData <= 1'b0;
            12'hbe6: oData <= 1'b0;
            12'hbe7: oData <= 1'b0;
            12'hbe8: oData <= 1'b0;
            12'hbe9: oData <= 1'b0;
            12'hbea: oData <= 1'b0;
            12'hbeb: oData <= 1'b0;
            12'hbec: oData <= 1'b0;
            12'hbed: oData <= 1'b0;
            12'hbee: oData <= 1'b0;
            12'hbef: oData <= 1'b0;
            12'hbf0: oData <= 1'b0;
            12'hbf1: oData <= 1'b0;
            12'hbf2: oData <= 1'b0;
            12'hbf3: oData <= 1'b0;
            12'hbf4: oData <= 1'b0;
            12'hbf5: oData <= 1'b0;
            12'hbf6: oData <= 1'b0;
            12'hbf7: oData <= 1'b0;
            12'hbf8: oData <= 1'b0;
            12'hbf9: oData <= 1'b0;
            12'hbfa: oData <= 1'b0;
            12'hbfb: oData <= 1'b0;
            12'hbfc: oData <= 1'b0;
            12'hbfd: oData <= 1'b0;
            12'hbfe: oData <= 1'b0;
            12'hbff: oData <= 1'b0;
            12'hc00: oData <= 1'b1;
            12'hc01: oData <= 1'b1;
            12'hc02: oData <= 1'b1;
            12'hc03: oData <= 1'b1;
            12'hc04: oData <= 1'b1;
            12'hc05: oData <= 1'b1;
            12'hc06: oData <= 1'b1;
            12'hc07: oData <= 1'b1;
            12'hc08: oData <= 1'b1;
            12'hc09: oData <= 1'b1;
            12'hc0a: oData <= 1'b1;
            12'hc0b: oData <= 1'b1;
            12'hc0c: oData <= 1'b1;
            12'hc0d: oData <= 1'b0;
            12'hc0e: oData <= 1'b0;
            12'hc0f: oData <= 1'b0;
            12'hc10: oData <= 1'b1;
            12'hc11: oData <= 1'b1;
            12'hc12: oData <= 1'b1;
            12'hc13: oData <= 1'b1;
            12'hc14: oData <= 1'b1;
            12'hc15: oData <= 1'b1;
            12'hc16: oData <= 1'b1;
            12'hc17: oData <= 1'b1;
            12'hc18: oData <= 1'b1;
            12'hc19: oData <= 1'b1;
            12'hc1a: oData <= 1'b1;
            12'hc1b: oData <= 1'b1;
            12'hc1c: oData <= 1'b1;
            12'hc1d: oData <= 1'b0;
            12'hc1e: oData <= 1'b0;
            12'hc1f: oData <= 1'b0;
            12'hc20: oData <= 1'b1;
            12'hc21: oData <= 1'b1;
            12'hc22: oData <= 1'b1;
            12'hc23: oData <= 1'b1;
            12'hc24: oData <= 1'b1;
            12'hc25: oData <= 1'b1;
            12'hc26: oData <= 1'b1;
            12'hc27: oData <= 1'b1;
            12'hc28: oData <= 1'b1;
            12'hc29: oData <= 1'b1;
            12'hc2a: oData <= 1'b1;
            12'hc2b: oData <= 1'b1;
            12'hc2c: oData <= 1'b1;
            12'hc2d: oData <= 1'b0;
            12'hc2e: oData <= 1'b0;
            12'hc2f: oData <= 1'b0;
            12'hc30: oData <= 1'b1;
            12'hc31: oData <= 1'b1;
            12'hc32: oData <= 1'b1;
            12'hc33: oData <= 1'b1;
            12'hc34: oData <= 1'b1;
            12'hc35: oData <= 1'b1;
            12'hc36: oData <= 1'b1;
            12'hc37: oData <= 1'b1;
            12'hc38: oData <= 1'b1;
            12'hc39: oData <= 1'b1;
            12'hc3a: oData <= 1'b1;
            12'hc3b: oData <= 1'b1;
            12'hc3c: oData <= 1'b1;
            12'hc3d: oData <= 1'b0;
            12'hc3e: oData <= 1'b0;
            12'hc3f: oData <= 1'b0;
            12'hc40: oData <= 1'b1;
            12'hc41: oData <= 1'b1;
            12'hc42: oData <= 1'b1;
            12'hc43: oData <= 1'b1;
            12'hc44: oData <= 1'b1;
            12'hc45: oData <= 1'b1;
            12'hc46: oData <= 1'b1;
            12'hc47: oData <= 1'b1;
            12'hc48: oData <= 1'b1;
            12'hc49: oData <= 1'b1;
            12'hc4a: oData <= 1'b1;
            12'hc4b: oData <= 1'b1;
            12'hc4c: oData <= 1'b0;
            12'hc4d: oData <= 1'b0;
            12'hc4e: oData <= 1'b0;
            12'hc4f: oData <= 1'b0;
            12'hc50: oData <= 1'b1;
            12'hc51: oData <= 1'b1;
            12'hc52: oData <= 1'b1;
            12'hc53: oData <= 1'b1;
            12'hc54: oData <= 1'b1;
            12'hc55: oData <= 1'b1;
            12'hc56: oData <= 1'b1;
            12'hc57: oData <= 1'b1;
            12'hc58: oData <= 1'b1;
            12'hc59: oData <= 1'b1;
            12'hc5a: oData <= 1'b1;
            12'hc5b: oData <= 1'b1;
            12'hc5c: oData <= 1'b0;
            12'hc5d: oData <= 1'b0;
            12'hc5e: oData <= 1'b0;
            12'hc5f: oData <= 1'b0;
            12'hc60: oData <= 1'b1;
            12'hc61: oData <= 1'b1;
            12'hc62: oData <= 1'b1;
            12'hc63: oData <= 1'b1;
            12'hc64: oData <= 1'b1;
            12'hc65: oData <= 1'b1;
            12'hc66: oData <= 1'b1;
            12'hc67: oData <= 1'b1;
            12'hc68: oData <= 1'b1;
            12'hc69: oData <= 1'b1;
            12'hc6a: oData <= 1'b1;
            12'hc6b: oData <= 1'b1;
            12'hc6c: oData <= 1'b0;
            12'hc6d: oData <= 1'b0;
            12'hc6e: oData <= 1'b0;
            12'hc6f: oData <= 1'b0;
            12'hc70: oData <= 1'b1;
            12'hc71: oData <= 1'b1;
            12'hc72: oData <= 1'b1;
            12'hc73: oData <= 1'b1;
            12'hc74: oData <= 1'b1;
            12'hc75: oData <= 1'b1;
            12'hc76: oData <= 1'b1;
            12'hc77: oData <= 1'b1;
            12'hc78: oData <= 1'b1;
            12'hc79: oData <= 1'b1;
            12'hc7a: oData <= 1'b1;
            12'hc7b: oData <= 1'b0;
            12'hc7c: oData <= 1'b0;
            12'hc7d: oData <= 1'b0;
            12'hc7e: oData <= 1'b0;
            12'hc7f: oData <= 1'b0;
            12'hc80: oData <= 1'b1;
            12'hc81: oData <= 1'b1;
            12'hc82: oData <= 1'b1;
            12'hc83: oData <= 1'b1;
            12'hc84: oData <= 1'b1;
            12'hc85: oData <= 1'b1;
            12'hc86: oData <= 1'b1;
            12'hc87: oData <= 1'b1;
            12'hc88: oData <= 1'b1;
            12'hc89: oData <= 1'b1;
            12'hc8a: oData <= 1'b1;
            12'hc8b: oData <= 1'b0;
            12'hc8c: oData <= 1'b0;
            12'hc8d: oData <= 1'b0;
            12'hc8e: oData <= 1'b0;
            12'hc8f: oData <= 1'b0;
            12'hc90: oData <= 1'b1;
            12'hc91: oData <= 1'b1;
            12'hc92: oData <= 1'b1;
            12'hc93: oData <= 1'b1;
            12'hc94: oData <= 1'b1;
            12'hc95: oData <= 1'b1;
            12'hc96: oData <= 1'b1;
            12'hc97: oData <= 1'b1;
            12'hc98: oData <= 1'b1;
            12'hc99: oData <= 1'b1;
            12'hc9a: oData <= 1'b0;
            12'hc9b: oData <= 1'b0;
            12'hc9c: oData <= 1'b0;
            12'hc9d: oData <= 1'b0;
            12'hc9e: oData <= 1'b0;
            12'hc9f: oData <= 1'b0;
            12'hca0: oData <= 1'b1;
            12'hca1: oData <= 1'b1;
            12'hca2: oData <= 1'b1;
            12'hca3: oData <= 1'b1;
            12'hca4: oData <= 1'b1;
            12'hca5: oData <= 1'b1;
            12'hca6: oData <= 1'b1;
            12'hca7: oData <= 1'b1;
            12'hca8: oData <= 1'b1;
            12'hca9: oData <= 1'b0;
            12'hcaa: oData <= 1'b0;
            12'hcab: oData <= 1'b0;
            12'hcac: oData <= 1'b0;
            12'hcad: oData <= 1'b0;
            12'hcae: oData <= 1'b0;
            12'hcaf: oData <= 1'b0;
            12'hcb0: oData <= 1'b1;
            12'hcb1: oData <= 1'b1;
            12'hcb2: oData <= 1'b1;
            12'hcb3: oData <= 1'b1;
            12'hcb4: oData <= 1'b1;
            12'hcb5: oData <= 1'b1;
            12'hcb6: oData <= 1'b1;
            12'hcb7: oData <= 1'b0;
            12'hcb8: oData <= 1'b0;
            12'hcb9: oData <= 1'b0;
            12'hcba: oData <= 1'b0;
            12'hcbb: oData <= 1'b0;
            12'hcbc: oData <= 1'b0;
            12'hcbd: oData <= 1'b0;
            12'hcbe: oData <= 1'b0;
            12'hcbf: oData <= 1'b0;
            12'hcc0: oData <= 1'b1;
            12'hcc1: oData <= 1'b1;
            12'hcc2: oData <= 1'b1;
            12'hcc3: oData <= 1'b1;
            12'hcc4: oData <= 1'b0;
            12'hcc5: oData <= 1'b0;
            12'hcc6: oData <= 1'b0;
            12'hcc7: oData <= 1'b0;
            12'hcc8: oData <= 1'b0;
            12'hcc9: oData <= 1'b0;
            12'hcca: oData <= 1'b0;
            12'hccb: oData <= 1'b0;
            12'hccc: oData <= 1'b0;
            12'hccd: oData <= 1'b0;
            12'hcce: oData <= 1'b0;
            12'hccf: oData <= 1'b0;
            12'hcd0: oData <= 1'b0;
            12'hcd1: oData <= 1'b0;
            12'hcd2: oData <= 1'b0;
            12'hcd3: oData <= 1'b0;
            12'hcd4: oData <= 1'b0;
            12'hcd5: oData <= 1'b0;
            12'hcd6: oData <= 1'b0;
            12'hcd7: oData <= 1'b0;
            12'hcd8: oData <= 1'b0;
            12'hcd9: oData <= 1'b0;
            12'hcda: oData <= 1'b0;
            12'hcdb: oData <= 1'b0;
            12'hcdc: oData <= 1'b0;
            12'hcdd: oData <= 1'b0;
            12'hcde: oData <= 1'b0;
            12'hcdf: oData <= 1'b0;
            12'hce0: oData <= 1'b0;
            12'hce1: oData <= 1'b0;
            12'hce2: oData <= 1'b0;
            12'hce3: oData <= 1'b0;
            12'hce4: oData <= 1'b0;
            12'hce5: oData <= 1'b0;
            12'hce6: oData <= 1'b0;
            12'hce7: oData <= 1'b0;
            12'hce8: oData <= 1'b0;
            12'hce9: oData <= 1'b0;
            12'hcea: oData <= 1'b0;
            12'hceb: oData <= 1'b0;
            12'hcec: oData <= 1'b0;
            12'hced: oData <= 1'b0;
            12'hcee: oData <= 1'b0;
            12'hcef: oData <= 1'b0;
            12'hcf0: oData <= 1'b0;
            12'hcf1: oData <= 1'b0;
            12'hcf2: oData <= 1'b0;
            12'hcf3: oData <= 1'b0;
            12'hcf4: oData <= 1'b0;
            12'hcf5: oData <= 1'b0;
            12'hcf6: oData <= 1'b0;
            12'hcf7: oData <= 1'b0;
            12'hcf8: oData <= 1'b0;
            12'hcf9: oData <= 1'b0;
            12'hcfa: oData <= 1'b0;
            12'hcfb: oData <= 1'b0;
            12'hcfc: oData <= 1'b0;
            12'hcfd: oData <= 1'b0;
            12'hcfe: oData <= 1'b0;
            12'hcff: oData <= 1'b0;
            12'hd00: oData <= 1'b1;
            12'hd01: oData <= 1'b1;
            12'hd02: oData <= 1'b1;
            12'hd03: oData <= 1'b1;
            12'hd04: oData <= 1'b1;
            12'hd05: oData <= 1'b1;
            12'hd06: oData <= 1'b1;
            12'hd07: oData <= 1'b1;
            12'hd08: oData <= 1'b1;
            12'hd09: oData <= 1'b1;
            12'hd0a: oData <= 1'b1;
            12'hd0b: oData <= 1'b1;
            12'hd0c: oData <= 1'b1;
            12'hd0d: oData <= 1'b1;
            12'hd0e: oData <= 1'b0;
            12'hd0f: oData <= 1'b0;
            12'hd10: oData <= 1'b1;
            12'hd11: oData <= 1'b1;
            12'hd12: oData <= 1'b1;
            12'hd13: oData <= 1'b1;
            12'hd14: oData <= 1'b1;
            12'hd15: oData <= 1'b1;
            12'hd16: oData <= 1'b1;
            12'hd17: oData <= 1'b1;
            12'hd18: oData <= 1'b1;
            12'hd19: oData <= 1'b1;
            12'hd1a: oData <= 1'b1;
            12'hd1b: oData <= 1'b1;
            12'hd1c: oData <= 1'b1;
            12'hd1d: oData <= 1'b1;
            12'hd1e: oData <= 1'b0;
            12'hd1f: oData <= 1'b0;
            12'hd20: oData <= 1'b1;
            12'hd21: oData <= 1'b1;
            12'hd22: oData <= 1'b1;
            12'hd23: oData <= 1'b1;
            12'hd24: oData <= 1'b1;
            12'hd25: oData <= 1'b1;
            12'hd26: oData <= 1'b1;
            12'hd27: oData <= 1'b1;
            12'hd28: oData <= 1'b1;
            12'hd29: oData <= 1'b1;
            12'hd2a: oData <= 1'b1;
            12'hd2b: oData <= 1'b1;
            12'hd2c: oData <= 1'b1;
            12'hd2d: oData <= 1'b1;
            12'hd2e: oData <= 1'b0;
            12'hd2f: oData <= 1'b0;
            12'hd30: oData <= 1'b1;
            12'hd31: oData <= 1'b1;
            12'hd32: oData <= 1'b1;
            12'hd33: oData <= 1'b1;
            12'hd34: oData <= 1'b1;
            12'hd35: oData <= 1'b1;
            12'hd36: oData <= 1'b1;
            12'hd37: oData <= 1'b1;
            12'hd38: oData <= 1'b1;
            12'hd39: oData <= 1'b1;
            12'hd3a: oData <= 1'b1;
            12'hd3b: oData <= 1'b1;
            12'hd3c: oData <= 1'b1;
            12'hd3d: oData <= 1'b1;
            12'hd3e: oData <= 1'b0;
            12'hd3f: oData <= 1'b0;
            12'hd40: oData <= 1'b1;
            12'hd41: oData <= 1'b1;
            12'hd42: oData <= 1'b1;
            12'hd43: oData <= 1'b1;
            12'hd44: oData <= 1'b1;
            12'hd45: oData <= 1'b1;
            12'hd46: oData <= 1'b1;
            12'hd47: oData <= 1'b1;
            12'hd48: oData <= 1'b1;
            12'hd49: oData <= 1'b1;
            12'hd4a: oData <= 1'b1;
            12'hd4b: oData <= 1'b1;
            12'hd4c: oData <= 1'b1;
            12'hd4d: oData <= 1'b0;
            12'hd4e: oData <= 1'b0;
            12'hd4f: oData <= 1'b0;
            12'hd50: oData <= 1'b1;
            12'hd51: oData <= 1'b1;
            12'hd52: oData <= 1'b1;
            12'hd53: oData <= 1'b1;
            12'hd54: oData <= 1'b1;
            12'hd55: oData <= 1'b1;
            12'hd56: oData <= 1'b1;
            12'hd57: oData <= 1'b1;
            12'hd58: oData <= 1'b1;
            12'hd59: oData <= 1'b1;
            12'hd5a: oData <= 1'b1;
            12'hd5b: oData <= 1'b1;
            12'hd5c: oData <= 1'b1;
            12'hd5d: oData <= 1'b0;
            12'hd5e: oData <= 1'b0;
            12'hd5f: oData <= 1'b0;
            12'hd60: oData <= 1'b1;
            12'hd61: oData <= 1'b1;
            12'hd62: oData <= 1'b1;
            12'hd63: oData <= 1'b1;
            12'hd64: oData <= 1'b1;
            12'hd65: oData <= 1'b1;
            12'hd66: oData <= 1'b1;
            12'hd67: oData <= 1'b1;
            12'hd68: oData <= 1'b1;
            12'hd69: oData <= 1'b1;
            12'hd6a: oData <= 1'b1;
            12'hd6b: oData <= 1'b1;
            12'hd6c: oData <= 1'b1;
            12'hd6d: oData <= 1'b0;
            12'hd6e: oData <= 1'b0;
            12'hd6f: oData <= 1'b0;
            12'hd70: oData <= 1'b1;
            12'hd71: oData <= 1'b1;
            12'hd72: oData <= 1'b1;
            12'hd73: oData <= 1'b1;
            12'hd74: oData <= 1'b1;
            12'hd75: oData <= 1'b1;
            12'hd76: oData <= 1'b1;
            12'hd77: oData <= 1'b1;
            12'hd78: oData <= 1'b1;
            12'hd79: oData <= 1'b1;
            12'hd7a: oData <= 1'b1;
            12'hd7b: oData <= 1'b1;
            12'hd7c: oData <= 1'b0;
            12'hd7d: oData <= 1'b0;
            12'hd7e: oData <= 1'b0;
            12'hd7f: oData <= 1'b0;
            12'hd80: oData <= 1'b1;
            12'hd81: oData <= 1'b1;
            12'hd82: oData <= 1'b1;
            12'hd83: oData <= 1'b1;
            12'hd84: oData <= 1'b1;
            12'hd85: oData <= 1'b1;
            12'hd86: oData <= 1'b1;
            12'hd87: oData <= 1'b1;
            12'hd88: oData <= 1'b1;
            12'hd89: oData <= 1'b1;
            12'hd8a: oData <= 1'b1;
            12'hd8b: oData <= 1'b1;
            12'hd8c: oData <= 1'b0;
            12'hd8d: oData <= 1'b0;
            12'hd8e: oData <= 1'b0;
            12'hd8f: oData <= 1'b0;
            12'hd90: oData <= 1'b1;
            12'hd91: oData <= 1'b1;
            12'hd92: oData <= 1'b1;
            12'hd93: oData <= 1'b1;
            12'hd94: oData <= 1'b1;
            12'hd95: oData <= 1'b1;
            12'hd96: oData <= 1'b1;
            12'hd97: oData <= 1'b1;
            12'hd98: oData <= 1'b1;
            12'hd99: oData <= 1'b1;
            12'hd9a: oData <= 1'b1;
            12'hd9b: oData <= 1'b0;
            12'hd9c: oData <= 1'b0;
            12'hd9d: oData <= 1'b0;
            12'hd9e: oData <= 1'b0;
            12'hd9f: oData <= 1'b0;
            12'hda0: oData <= 1'b1;
            12'hda1: oData <= 1'b1;
            12'hda2: oData <= 1'b1;
            12'hda3: oData <= 1'b1;
            12'hda4: oData <= 1'b1;
            12'hda5: oData <= 1'b1;
            12'hda6: oData <= 1'b1;
            12'hda7: oData <= 1'b1;
            12'hda8: oData <= 1'b1;
            12'hda9: oData <= 1'b1;
            12'hdaa: oData <= 1'b0;
            12'hdab: oData <= 1'b0;
            12'hdac: oData <= 1'b0;
            12'hdad: oData <= 1'b0;
            12'hdae: oData <= 1'b0;
            12'hdaf: oData <= 1'b0;
            12'hdb0: oData <= 1'b1;
            12'hdb1: oData <= 1'b1;
            12'hdb2: oData <= 1'b1;
            12'hdb3: oData <= 1'b1;
            12'hdb4: oData <= 1'b1;
            12'hdb5: oData <= 1'b1;
            12'hdb6: oData <= 1'b1;
            12'hdb7: oData <= 1'b1;
            12'hdb8: oData <= 1'b1;
            12'hdb9: oData <= 1'b0;
            12'hdba: oData <= 1'b0;
            12'hdbb: oData <= 1'b0;
            12'hdbc: oData <= 1'b0;
            12'hdbd: oData <= 1'b0;
            12'hdbe: oData <= 1'b0;
            12'hdbf: oData <= 1'b0;
            12'hdc0: oData <= 1'b1;
            12'hdc1: oData <= 1'b1;
            12'hdc2: oData <= 1'b1;
            12'hdc3: oData <= 1'b1;
            12'hdc4: oData <= 1'b1;
            12'hdc5: oData <= 1'b1;
            12'hdc6: oData <= 1'b1;
            12'hdc7: oData <= 1'b0;
            12'hdc8: oData <= 1'b0;
            12'hdc9: oData <= 1'b0;
            12'hdca: oData <= 1'b0;
            12'hdcb: oData <= 1'b0;
            12'hdcc: oData <= 1'b0;
            12'hdcd: oData <= 1'b0;
            12'hdce: oData <= 1'b0;
            12'hdcf: oData <= 1'b0;
            12'hdd0: oData <= 1'b1;
            12'hdd1: oData <= 1'b1;
            12'hdd2: oData <= 1'b1;
            12'hdd3: oData <= 1'b1;
            12'hdd4: oData <= 1'b0;
            12'hdd5: oData <= 1'b0;
            12'hdd6: oData <= 1'b0;
            12'hdd7: oData <= 1'b0;
            12'hdd8: oData <= 1'b0;
            12'hdd9: oData <= 1'b0;
            12'hdda: oData <= 1'b0;
            12'hddb: oData <= 1'b0;
            12'hddc: oData <= 1'b0;
            12'hddd: oData <= 1'b0;
            12'hdde: oData <= 1'b0;
            12'hddf: oData <= 1'b0;
            12'hde0: oData <= 1'b0;
            12'hde1: oData <= 1'b0;
            12'hde2: oData <= 1'b0;
            12'hde3: oData <= 1'b0;
            12'hde4: oData <= 1'b0;
            12'hde5: oData <= 1'b0;
            12'hde6: oData <= 1'b0;
            12'hde7: oData <= 1'b0;
            12'hde8: oData <= 1'b0;
            12'hde9: oData <= 1'b0;
            12'hdea: oData <= 1'b0;
            12'hdeb: oData <= 1'b0;
            12'hdec: oData <= 1'b0;
            12'hded: oData <= 1'b0;
            12'hdee: oData <= 1'b0;
            12'hdef: oData <= 1'b0;
            12'hdf0: oData <= 1'b0;
            12'hdf1: oData <= 1'b0;
            12'hdf2: oData <= 1'b0;
            12'hdf3: oData <= 1'b0;
            12'hdf4: oData <= 1'b0;
            12'hdf5: oData <= 1'b0;
            12'hdf6: oData <= 1'b0;
            12'hdf7: oData <= 1'b0;
            12'hdf8: oData <= 1'b0;
            12'hdf9: oData <= 1'b0;
            12'hdfa: oData <= 1'b0;
            12'hdfb: oData <= 1'b0;
            12'hdfc: oData <= 1'b0;
            12'hdfd: oData <= 1'b0;
            12'hdfe: oData <= 1'b0;
            12'hdff: oData <= 1'b0;
            12'he00: oData <= 1'b1;
            12'he01: oData <= 1'b1;
            12'he02: oData <= 1'b1;
            12'he03: oData <= 1'b1;
            12'he04: oData <= 1'b1;
            12'he05: oData <= 1'b1;
            12'he06: oData <= 1'b1;
            12'he07: oData <= 1'b1;
            12'he08: oData <= 1'b1;
            12'he09: oData <= 1'b1;
            12'he0a: oData <= 1'b1;
            12'he0b: oData <= 1'b1;
            12'he0c: oData <= 1'b1;
            12'he0d: oData <= 1'b1;
            12'he0e: oData <= 1'b1;
            12'he0f: oData <= 1'b0;
            12'he10: oData <= 1'b1;
            12'he11: oData <= 1'b1;
            12'he12: oData <= 1'b1;
            12'he13: oData <= 1'b1;
            12'he14: oData <= 1'b1;
            12'he15: oData <= 1'b1;
            12'he16: oData <= 1'b1;
            12'he17: oData <= 1'b1;
            12'he18: oData <= 1'b1;
            12'he19: oData <= 1'b1;
            12'he1a: oData <= 1'b1;
            12'he1b: oData <= 1'b1;
            12'he1c: oData <= 1'b1;
            12'he1d: oData <= 1'b1;
            12'he1e: oData <= 1'b1;
            12'he1f: oData <= 1'b0;
            12'he20: oData <= 1'b1;
            12'he21: oData <= 1'b1;
            12'he22: oData <= 1'b1;
            12'he23: oData <= 1'b1;
            12'he24: oData <= 1'b1;
            12'he25: oData <= 1'b1;
            12'he26: oData <= 1'b1;
            12'he27: oData <= 1'b1;
            12'he28: oData <= 1'b1;
            12'he29: oData <= 1'b1;
            12'he2a: oData <= 1'b1;
            12'he2b: oData <= 1'b1;
            12'he2c: oData <= 1'b1;
            12'he2d: oData <= 1'b1;
            12'he2e: oData <= 1'b1;
            12'he2f: oData <= 1'b0;
            12'he30: oData <= 1'b1;
            12'he31: oData <= 1'b1;
            12'he32: oData <= 1'b1;
            12'he33: oData <= 1'b1;
            12'he34: oData <= 1'b1;
            12'he35: oData <= 1'b1;
            12'he36: oData <= 1'b1;
            12'he37: oData <= 1'b1;
            12'he38: oData <= 1'b1;
            12'he39: oData <= 1'b1;
            12'he3a: oData <= 1'b1;
            12'he3b: oData <= 1'b1;
            12'he3c: oData <= 1'b1;
            12'he3d: oData <= 1'b1;
            12'he3e: oData <= 1'b1;
            12'he3f: oData <= 1'b0;
            12'he40: oData <= 1'b1;
            12'he41: oData <= 1'b1;
            12'he42: oData <= 1'b1;
            12'he43: oData <= 1'b1;
            12'he44: oData <= 1'b1;
            12'he45: oData <= 1'b1;
            12'he46: oData <= 1'b1;
            12'he47: oData <= 1'b1;
            12'he48: oData <= 1'b1;
            12'he49: oData <= 1'b1;
            12'he4a: oData <= 1'b1;
            12'he4b: oData <= 1'b1;
            12'he4c: oData <= 1'b1;
            12'he4d: oData <= 1'b1;
            12'he4e: oData <= 1'b0;
            12'he4f: oData <= 1'b0;
            12'he50: oData <= 1'b1;
            12'he51: oData <= 1'b1;
            12'he52: oData <= 1'b1;
            12'he53: oData <= 1'b1;
            12'he54: oData <= 1'b1;
            12'he55: oData <= 1'b1;
            12'he56: oData <= 1'b1;
            12'he57: oData <= 1'b1;
            12'he58: oData <= 1'b1;
            12'he59: oData <= 1'b1;
            12'he5a: oData <= 1'b1;
            12'he5b: oData <= 1'b1;
            12'he5c: oData <= 1'b1;
            12'he5d: oData <= 1'b1;
            12'he5e: oData <= 1'b0;
            12'he5f: oData <= 1'b0;
            12'he60: oData <= 1'b1;
            12'he61: oData <= 1'b1;
            12'he62: oData <= 1'b1;
            12'he63: oData <= 1'b1;
            12'he64: oData <= 1'b1;
            12'he65: oData <= 1'b1;
            12'he66: oData <= 1'b1;
            12'he67: oData <= 1'b1;
            12'he68: oData <= 1'b1;
            12'he69: oData <= 1'b1;
            12'he6a: oData <= 1'b1;
            12'he6b: oData <= 1'b1;
            12'he6c: oData <= 1'b1;
            12'he6d: oData <= 1'b1;
            12'he6e: oData <= 1'b0;
            12'he6f: oData <= 1'b0;
            12'he70: oData <= 1'b1;
            12'he71: oData <= 1'b1;
            12'he72: oData <= 1'b1;
            12'he73: oData <= 1'b1;
            12'he74: oData <= 1'b1;
            12'he75: oData <= 1'b1;
            12'he76: oData <= 1'b1;
            12'he77: oData <= 1'b1;
            12'he78: oData <= 1'b1;
            12'he79: oData <= 1'b1;
            12'he7a: oData <= 1'b1;
            12'he7b: oData <= 1'b1;
            12'he7c: oData <= 1'b1;
            12'he7d: oData <= 1'b0;
            12'he7e: oData <= 1'b0;
            12'he7f: oData <= 1'b0;
            12'he80: oData <= 1'b1;
            12'he81: oData <= 1'b1;
            12'he82: oData <= 1'b1;
            12'he83: oData <= 1'b1;
            12'he84: oData <= 1'b1;
            12'he85: oData <= 1'b1;
            12'he86: oData <= 1'b1;
            12'he87: oData <= 1'b1;
            12'he88: oData <= 1'b1;
            12'he89: oData <= 1'b1;
            12'he8a: oData <= 1'b1;
            12'he8b: oData <= 1'b1;
            12'he8c: oData <= 1'b1;
            12'he8d: oData <= 1'b0;
            12'he8e: oData <= 1'b0;
            12'he8f: oData <= 1'b0;
            12'he90: oData <= 1'b1;
            12'he91: oData <= 1'b1;
            12'he92: oData <= 1'b1;
            12'he93: oData <= 1'b1;
            12'he94: oData <= 1'b1;
            12'he95: oData <= 1'b1;
            12'he96: oData <= 1'b1;
            12'he97: oData <= 1'b1;
            12'he98: oData <= 1'b1;
            12'he99: oData <= 1'b1;
            12'he9a: oData <= 1'b1;
            12'he9b: oData <= 1'b1;
            12'he9c: oData <= 1'b0;
            12'he9d: oData <= 1'b0;
            12'he9e: oData <= 1'b0;
            12'he9f: oData <= 1'b0;
            12'hea0: oData <= 1'b1;
            12'hea1: oData <= 1'b1;
            12'hea2: oData <= 1'b1;
            12'hea3: oData <= 1'b1;
            12'hea4: oData <= 1'b1;
            12'hea5: oData <= 1'b1;
            12'hea6: oData <= 1'b1;
            12'hea7: oData <= 1'b1;
            12'hea8: oData <= 1'b1;
            12'hea9: oData <= 1'b1;
            12'heaa: oData <= 1'b1;
            12'heab: oData <= 1'b0;
            12'heac: oData <= 1'b0;
            12'head: oData <= 1'b0;
            12'heae: oData <= 1'b0;
            12'heaf: oData <= 1'b0;
            12'heb0: oData <= 1'b1;
            12'heb1: oData <= 1'b1;
            12'heb2: oData <= 1'b1;
            12'heb3: oData <= 1'b1;
            12'heb4: oData <= 1'b1;
            12'heb5: oData <= 1'b1;
            12'heb6: oData <= 1'b1;
            12'heb7: oData <= 1'b1;
            12'heb8: oData <= 1'b1;
            12'heb9: oData <= 1'b1;
            12'heba: oData <= 1'b0;
            12'hebb: oData <= 1'b0;
            12'hebc: oData <= 1'b0;
            12'hebd: oData <= 1'b0;
            12'hebe: oData <= 1'b0;
            12'hebf: oData <= 1'b0;
            12'hec0: oData <= 1'b1;
            12'hec1: oData <= 1'b1;
            12'hec2: oData <= 1'b1;
            12'hec3: oData <= 1'b1;
            12'hec4: oData <= 1'b1;
            12'hec5: oData <= 1'b1;
            12'hec6: oData <= 1'b1;
            12'hec7: oData <= 1'b1;
            12'hec8: oData <= 1'b1;
            12'hec9: oData <= 1'b0;
            12'heca: oData <= 1'b0;
            12'hecb: oData <= 1'b0;
            12'hecc: oData <= 1'b0;
            12'hecd: oData <= 1'b0;
            12'hece: oData <= 1'b0;
            12'hecf: oData <= 1'b0;
            12'hed0: oData <= 1'b1;
            12'hed1: oData <= 1'b1;
            12'hed2: oData <= 1'b1;
            12'hed3: oData <= 1'b1;
            12'hed4: oData <= 1'b1;
            12'hed5: oData <= 1'b1;
            12'hed6: oData <= 1'b1;
            12'hed7: oData <= 1'b0;
            12'hed8: oData <= 1'b0;
            12'hed9: oData <= 1'b0;
            12'heda: oData <= 1'b0;
            12'hedb: oData <= 1'b0;
            12'hedc: oData <= 1'b0;
            12'hedd: oData <= 1'b0;
            12'hede: oData <= 1'b0;
            12'hedf: oData <= 1'b0;
            12'hee0: oData <= 1'b1;
            12'hee1: oData <= 1'b1;
            12'hee2: oData <= 1'b1;
            12'hee3: oData <= 1'b1;
            12'hee4: oData <= 1'b0;
            12'hee5: oData <= 1'b0;
            12'hee6: oData <= 1'b0;
            12'hee7: oData <= 1'b0;
            12'hee8: oData <= 1'b0;
            12'hee9: oData <= 1'b0;
            12'heea: oData <= 1'b0;
            12'heeb: oData <= 1'b0;
            12'heec: oData <= 1'b0;
            12'heed: oData <= 1'b0;
            12'heee: oData <= 1'b0;
            12'heef: oData <= 1'b0;
            12'hef0: oData <= 1'b0;
            12'hef1: oData <= 1'b0;
            12'hef2: oData <= 1'b0;
            12'hef3: oData <= 1'b0;
            12'hef4: oData <= 1'b0;
            12'hef5: oData <= 1'b0;
            12'hef6: oData <= 1'b0;
            12'hef7: oData <= 1'b0;
            12'hef8: oData <= 1'b0;
            12'hef9: oData <= 1'b0;
            12'hefa: oData <= 1'b0;
            12'hefb: oData <= 1'b0;
            12'hefc: oData <= 1'b0;
            12'hefd: oData <= 1'b0;
            12'hefe: oData <= 1'b0;
            12'heff: oData <= 1'b0;
            12'hf00: oData <= 1'b1;
            12'hf01: oData <= 1'b1;
            12'hf02: oData <= 1'b1;
            12'hf03: oData <= 1'b1;
            12'hf04: oData <= 1'b1;
            12'hf05: oData <= 1'b1;
            12'hf06: oData <= 1'b1;
            12'hf07: oData <= 1'b1;
            12'hf08: oData <= 1'b1;
            12'hf09: oData <= 1'b1;
            12'hf0a: oData <= 1'b1;
            12'hf0b: oData <= 1'b1;
            12'hf0c: oData <= 1'b1;
            12'hf0d: oData <= 1'b1;
            12'hf0e: oData <= 1'b1;
            12'hf0f: oData <= 1'b1;
            12'hf10: oData <= 1'b1;
            12'hf11: oData <= 1'b1;
            12'hf12: oData <= 1'b1;
            12'hf13: oData <= 1'b1;
            12'hf14: oData <= 1'b1;
            12'hf15: oData <= 1'b1;
            12'hf16: oData <= 1'b1;
            12'hf17: oData <= 1'b1;
            12'hf18: oData <= 1'b1;
            12'hf19: oData <= 1'b1;
            12'hf1a: oData <= 1'b1;
            12'hf1b: oData <= 1'b1;
            12'hf1c: oData <= 1'b1;
            12'hf1d: oData <= 1'b1;
            12'hf1e: oData <= 1'b1;
            12'hf1f: oData <= 1'b1;
            12'hf20: oData <= 1'b1;
            12'hf21: oData <= 1'b1;
            12'hf22: oData <= 1'b1;
            12'hf23: oData <= 1'b1;
            12'hf24: oData <= 1'b1;
            12'hf25: oData <= 1'b1;
            12'hf26: oData <= 1'b1;
            12'hf27: oData <= 1'b1;
            12'hf28: oData <= 1'b1;
            12'hf29: oData <= 1'b1;
            12'hf2a: oData <= 1'b1;
            12'hf2b: oData <= 1'b1;
            12'hf2c: oData <= 1'b1;
            12'hf2d: oData <= 1'b1;
            12'hf2e: oData <= 1'b1;
            12'hf2f: oData <= 1'b1;
            12'hf30: oData <= 1'b1;
            12'hf31: oData <= 1'b1;
            12'hf32: oData <= 1'b1;
            12'hf33: oData <= 1'b1;
            12'hf34: oData <= 1'b1;
            12'hf35: oData <= 1'b1;
            12'hf36: oData <= 1'b1;
            12'hf37: oData <= 1'b1;
            12'hf38: oData <= 1'b1;
            12'hf39: oData <= 1'b1;
            12'hf3a: oData <= 1'b1;
            12'hf3b: oData <= 1'b1;
            12'hf3c: oData <= 1'b1;
            12'hf3d: oData <= 1'b1;
            12'hf3e: oData <= 1'b1;
            12'hf3f: oData <= 1'b1;
            12'hf40: oData <= 1'b1;
            12'hf41: oData <= 1'b1;
            12'hf42: oData <= 1'b1;
            12'hf43: oData <= 1'b1;
            12'hf44: oData <= 1'b1;
            12'hf45: oData <= 1'b1;
            12'hf46: oData <= 1'b1;
            12'hf47: oData <= 1'b1;
            12'hf48: oData <= 1'b1;
            12'hf49: oData <= 1'b1;
            12'hf4a: oData <= 1'b1;
            12'hf4b: oData <= 1'b1;
            12'hf4c: oData <= 1'b1;
            12'hf4d: oData <= 1'b1;
            12'hf4e: oData <= 1'b1;
            12'hf4f: oData <= 1'b1;
            12'hf50: oData <= 1'b1;
            12'hf51: oData <= 1'b1;
            12'hf52: oData <= 1'b1;
            12'hf53: oData <= 1'b1;
            12'hf54: oData <= 1'b1;
            12'hf55: oData <= 1'b1;
            12'hf56: oData <= 1'b1;
            12'hf57: oData <= 1'b1;
            12'hf58: oData <= 1'b1;
            12'hf59: oData <= 1'b1;
            12'hf5a: oData <= 1'b1;
            12'hf5b: oData <= 1'b1;
            12'hf5c: oData <= 1'b1;
            12'hf5d: oData <= 1'b1;
            12'hf5e: oData <= 1'b1;
            12'hf5f: oData <= 1'b0;
            12'hf60: oData <= 1'b1;
            12'hf61: oData <= 1'b1;
            12'hf62: oData <= 1'b1;
            12'hf63: oData <= 1'b1;
            12'hf64: oData <= 1'b1;
            12'hf65: oData <= 1'b1;
            12'hf66: oData <= 1'b1;
            12'hf67: oData <= 1'b1;
            12'hf68: oData <= 1'b1;
            12'hf69: oData <= 1'b1;
            12'hf6a: oData <= 1'b1;
            12'hf6b: oData <= 1'b1;
            12'hf6c: oData <= 1'b1;
            12'hf6d: oData <= 1'b1;
            12'hf6e: oData <= 1'b1;
            12'hf6f: oData <= 1'b0;
            12'hf70: oData <= 1'b1;
            12'hf71: oData <= 1'b1;
            12'hf72: oData <= 1'b1;
            12'hf73: oData <= 1'b1;
            12'hf74: oData <= 1'b1;
            12'hf75: oData <= 1'b1;
            12'hf76: oData <= 1'b1;
            12'hf77: oData <= 1'b1;
            12'hf78: oData <= 1'b1;
            12'hf79: oData <= 1'b1;
            12'hf7a: oData <= 1'b1;
            12'hf7b: oData <= 1'b1;
            12'hf7c: oData <= 1'b1;
            12'hf7d: oData <= 1'b1;
            12'hf7e: oData <= 1'b0;
            12'hf7f: oData <= 1'b0;
            12'hf80: oData <= 1'b1;
            12'hf81: oData <= 1'b1;
            12'hf82: oData <= 1'b1;
            12'hf83: oData <= 1'b1;
            12'hf84: oData <= 1'b1;
            12'hf85: oData <= 1'b1;
            12'hf86: oData <= 1'b1;
            12'hf87: oData <= 1'b1;
            12'hf88: oData <= 1'b1;
            12'hf89: oData <= 1'b1;
            12'hf8a: oData <= 1'b1;
            12'hf8b: oData <= 1'b1;
            12'hf8c: oData <= 1'b1;
            12'hf8d: oData <= 1'b1;
            12'hf8e: oData <= 1'b0;
            12'hf8f: oData <= 1'b0;
            12'hf90: oData <= 1'b1;
            12'hf91: oData <= 1'b1;
            12'hf92: oData <= 1'b1;
            12'hf93: oData <= 1'b1;
            12'hf94: oData <= 1'b1;
            12'hf95: oData <= 1'b1;
            12'hf96: oData <= 1'b1;
            12'hf97: oData <= 1'b1;
            12'hf98: oData <= 1'b1;
            12'hf99: oData <= 1'b1;
            12'hf9a: oData <= 1'b1;
            12'hf9b: oData <= 1'b1;
            12'hf9c: oData <= 1'b1;
            12'hf9d: oData <= 1'b0;
            12'hf9e: oData <= 1'b0;
            12'hf9f: oData <= 1'b0;
            12'hfa0: oData <= 1'b1;
            12'hfa1: oData <= 1'b1;
            12'hfa2: oData <= 1'b1;
            12'hfa3: oData <= 1'b1;
            12'hfa4: oData <= 1'b1;
            12'hfa5: oData <= 1'b1;
            12'hfa6: oData <= 1'b1;
            12'hfa7: oData <= 1'b1;
            12'hfa8: oData <= 1'b1;
            12'hfa9: oData <= 1'b1;
            12'hfaa: oData <= 1'b1;
            12'hfab: oData <= 1'b1;
            12'hfac: oData <= 1'b0;
            12'hfad: oData <= 1'b0;
            12'hfae: oData <= 1'b0;
            12'hfaf: oData <= 1'b0;
            12'hfb0: oData <= 1'b1;
            12'hfb1: oData <= 1'b1;
            12'hfb2: oData <= 1'b1;
            12'hfb3: oData <= 1'b1;
            12'hfb4: oData <= 1'b1;
            12'hfb5: oData <= 1'b1;
            12'hfb6: oData <= 1'b1;
            12'hfb7: oData <= 1'b1;
            12'hfb8: oData <= 1'b1;
            12'hfb9: oData <= 1'b1;
            12'hfba: oData <= 1'b1;
            12'hfbb: oData <= 1'b0;
            12'hfbc: oData <= 1'b0;
            12'hfbd: oData <= 1'b0;
            12'hfbe: oData <= 1'b0;
            12'hfbf: oData <= 1'b0;
            12'hfc0: oData <= 1'b1;
            12'hfc1: oData <= 1'b1;
            12'hfc2: oData <= 1'b1;
            12'hfc3: oData <= 1'b1;
            12'hfc4: oData <= 1'b1;
            12'hfc5: oData <= 1'b1;
            12'hfc6: oData <= 1'b1;
            12'hfc7: oData <= 1'b1;
            12'hfc8: oData <= 1'b1;
            12'hfc9: oData <= 1'b1;
            12'hfca: oData <= 1'b0;
            12'hfcb: oData <= 1'b0;
            12'hfcc: oData <= 1'b0;
            12'hfcd: oData <= 1'b0;
            12'hfce: oData <= 1'b0;
            12'hfcf: oData <= 1'b0;
            12'hfd0: oData <= 1'b1;
            12'hfd1: oData <= 1'b1;
            12'hfd2: oData <= 1'b1;
            12'hfd3: oData <= 1'b1;
            12'hfd4: oData <= 1'b1;
            12'hfd5: oData <= 1'b1;
            12'hfd6: oData <= 1'b1;
            12'hfd7: oData <= 1'b1;
            12'hfd8: oData <= 1'b1;
            12'hfd9: oData <= 1'b0;
            12'hfda: oData <= 1'b0;
            12'hfdb: oData <= 1'b0;
            12'hfdc: oData <= 1'b0;
            12'hfdd: oData <= 1'b0;
            12'hfde: oData <= 1'b0;
            12'hfdf: oData <= 1'b0;
            12'hfe0: oData <= 1'b1;
            12'hfe1: oData <= 1'b1;
            12'hfe2: oData <= 1'b1;
            12'hfe3: oData <= 1'b1;
            12'hfe4: oData <= 1'b1;
            12'hfe5: oData <= 1'b1;
            12'hfe6: oData <= 1'b1;
            12'hfe7: oData <= 1'b0;
            12'hfe8: oData <= 1'b0;
            12'hfe9: oData <= 1'b0;
            12'hfea: oData <= 1'b0;
            12'hfeb: oData <= 1'b0;
            12'hfec: oData <= 1'b0;
            12'hfed: oData <= 1'b0;
            12'hfee: oData <= 1'b0;
            12'hfef: oData <= 1'b0;
            12'hff0: oData <= 1'b1;
            12'hff1: oData <= 1'b1;
            12'hff2: oData <= 1'b1;
            12'hff3: oData <= 1'b1;
            12'hff4: oData <= 1'b1;
            12'hff5: oData <= 1'b0;
            12'hff6: oData <= 1'b0;
            12'hff7: oData <= 1'b0;
            12'hff8: oData <= 1'b0;
            12'hff9: oData <= 1'b0;
            12'hffa: oData <= 1'b0;
            12'hffb: oData <= 1'b0;
            12'hffc: oData <= 1'b0;
            12'hffd: oData <= 1'b0;
            12'hffe: oData <= 1'b0;
            12'hfff: oData <= 1'b0;
        endcase
    end
endmodule
