// megafunction wizard: %LPM_DIVIDE%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_divide 

// ============================================================
// File Name: divider7stage.v
// Megafunction Name(s):
// 			lpm_divide
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.0 Build 178 04/27/2006 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2006 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module divider5stage (
	clken,
	clock,
	denom,
	numer,
	quotient,
	remain);
	
parameter BusWidth = 0;
parameter DecimalWidth = 0;

	input	  clken;
	input	  clock;
	input	[BusWidth-1:0]  denom;
	input	[BusWidth+DecimalWidth-1:0]  numer;
	output	[BusWidth+DecimalWidth-1:0]  quotient;
	output	[BusWidth-1:0]  remain;

	wire [BusWidth+DecimalWidth-1:0] sub_wire0;
	wire [BusWidth-1:0] sub_wire1;
	wire [BusWidth+DecimalWidth-1:0] quotient = sub_wire0[BusWidth+DecimalWidth-1:0];
	wire [BusWidth-1:0] remain = sub_wire1[BusWidth-1:0];

	lpm_divide	lpm_divide_component (
				.clken (clken),
				.denom (denom),
				.clock (clock),
				.numer (numer),
				.quotient (sub_wire0),
				.remain (sub_wire1),
				.aclr (1'b0));
	defparam
		lpm_divide_component.lpm_drepresentation = "SIGNED",
		lpm_divide_component.lpm_hint = "MAXIMIZE_SPEED=6,LPM_REMAINDERPOSITIVE=FALSE",
		lpm_divide_component.lpm_nrepresentation = "SIGNED",
		lpm_divide_component.lpm_pipeline = 5,
		lpm_divide_component.lpm_type = "LPM_DIVIDE",
		lpm_divide_component.lpm_widthd = BusWidth,
		lpm_divide_component.lpm_widthn = BusWidth+DecimalWidth;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "FALSE"
// Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "6"
// Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1"
// Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
// Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=6,LPM_REMAINDERPOSITIVE=FALSE"
// Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "5"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
// Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "24"
// Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "40"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT NODEFVAL clken
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: denom 0 0 24 0 INPUT NODEFVAL denom[23..0]
// Retrieval info: USED_PORT: numer 0 0 40 0 INPUT NODEFVAL numer[39..0]
// Retrieval info: USED_PORT: quotient 0 0 40 0 OUTPUT NODEFVAL quotient[39..0]
// Retrieval info: USED_PORT: remain 0 0 24 0 OUTPUT NODEFVAL remain[23..0]
// Retrieval info: CONNECT: @numer 0 0 40 0 numer 0 0 40 0
// Retrieval info: CONNECT: @denom 0 0 24 0 denom 0 0 24 0
// Retrieval info: CONNECT: quotient 0 0 40 0 @quotient 0 0 40 0
// Retrieval info: CONNECT: remain 0 0 24 0 @remain 0 0 24 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL divider.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider_bb.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL divider5stage_bb.v FALSE
